--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v
X"3B9A",
X"0188",
X"0311",
X"0499",
X"0620",
X"07A6",
X"092B",
X"0AAF",
X"0C31",
X"0DB1",
X"0F2F",
X"10AB",
X"1224",
X"139A",
X"150E",
X"167E",
X"17EA",
X"1953",
X"1AB8",
X"1C19",
X"1D76",
X"1ECE",
X"2021",
X"216F",
X"22B9",
X"23FC",
X"253B",
X"2673",
X"27A6",
X"28D2",
X"29F8",
X"2B18",
X"2C31",
X"2D43",
X"2E4F",
X"2F53",
X"3050",
X"3145",
X"3233",
X"3319",
X"33F7",
X"34CD",
X"359B",
X"3661",
X"371E",
X"37D3",
X"387F",
X"3923",
X"39BE",
X"3A4F",
X"3AD8",
X"3B58",
X"3BCF",
X"3C3C",
X"3CA0",
X"3CFB",
X"3D4C",
X"3D94",
X"3DD2",
X"3E07",
X"3E32",
X"3E54",
X"3E6C",
X"3E7B",
X"3E80",
X"3E7B",
X"3E6C",
X"3E54",
X"3E32",
X"3E07",
X"3DD2",
X"3D94",
X"3D4C",
X"3CFB",
X"3CA0",
X"3C3C",
X"3BCF",
X"3B58",
X"3AD8",
X"3A4F",
X"39BE",
X"3923",
X"387F",
X"37D3",
X"371E",
X"3661",
X"359B",
X"34CD",
X"33F7",
X"3319",
X"3233",
X"3145",
X"3050",
X"2F53",
X"2E4F",
X"2D43",
X"2C31",
X"2B18",
X"29F8",
X"28D2",
X"27A6",
X"2673",
X"253B",
X"23FC",
X"22B9",
X"216F",
X"2021",
X"1ECE",
X"1D76",
X"1C19",
X"1AB8",
X"1953",
X"17EA",
X"167E",
X"150E",
X"139A",
X"1224",
X"10AB",
X"0F2F",
X"0DB1",
X"0C31",
X"0AAF",
X"092B",
X"07A6",
X"0620",
X"0499",
X"0311",
X"0188",
X"0000",
X"FE78",
X"FCEF",
X"FB67",
X"F9E0",
X"F85A",
X"F6D5",
X"F551",
X"F3CF",
X"F24F",
X"F0D1",
X"EF55",
X"EDDC",
X"EC66",
X"EAF2",
X"E982",
X"E816",
X"E6AD",
X"E548",
X"E3E7",
X"E28A",
X"E132",
X"DFDF",
X"DE91",
X"DD47",
X"DC04",
X"DAC5",
X"D98D",
X"D85A",
X"D72E",
X"D608",
X"D4E8",
X"D3CF",
X"D2BD",
X"D1B1",
X"D0AD",
X"CFB0",
X"CEBB",
X"CDCD",
X"CCE7",
X"CC09",
X"CB33",
X"CA65",
X"C99F",
X"C8E2",
X"C82D",
X"C781",
X"C6DD",
X"C642",
X"C5B1",
X"C528",
X"C4A8",
X"C431",
X"C3C4",
X"C360",
X"C305",
X"C2B4",
X"C26C",
X"C22E",
X"C1F9",
X"C1CE",
X"C1AC",
X"C194",
X"C185",
X"C180",
X"C185",
X"C194",
X"C1AC",
X"C1CE",
X"C1F9",
X"C22E",
X"C26C",
X"C2B4",
X"C305",
X"C360",
X"C3C4",
X"C431",
X"C4A8",
X"C528",
X"C5B1",
X"C642",
X"C6DD",
X"C781",
X"C82D",
X"C8E2",
X"C99F",
X"CA65",
X"CB33",
X"CC09",
X"CCE7",
X"CDCD",
X"CEBB",
X"CFB0",
X"D0AD",
X"D1B1",
X"D2BD",
X"D3CF",
X"D4E8",
X"D608",
X"D72E",
X"D85A",
X"D98D",
X"DAC5",
X"DC04",
X"DD47",
X"DE91",
X"DFDF",
X"E132",
X"E28A",
X"E3E7",
X"E548",
X"E6AD",
X"E816",
X"E982",
X"EAF2",
X"EC66",
X"EDDC",
X"EF55",
X"F0D1",
X"F24F",
X"F3CF",
X"F551",
X"F6D5",
X"F85A",
X"F9E0",
X"FB67",
X"FCEF",
X"FE78"


 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;