library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity blue_car_44_22_object is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end blue_car_44_22_object;

architecture behav of blue_car_44_22_object is

constant object_X_size : integer := 44;
constant object_Y_size : integer := 22;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"2E", x"29", x"37", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"20", x"00", x"04", x"09", x"29", x"2E", x"2E", x"2E", x"2E", x"2E", x"2E", x"2E", x"2D", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"09", x"33", x"32", x"05", x"29", x"29", x"29", x"29", x"2E", x"2E", x"2E", x"2E", x"2E", x"2E", x"29", x"00", x"2D", x"00", x"00", x"00"),
(x"00", x"09", x"2D", x"2E", x"33", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"32", x"29", x"00", x"00", x"00"),
(x"29", x"33", x"37", x"37", x"3B", x"3B", x"3B", x"37", x"37", x"37", x"37", x"37", x"32", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"2E", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"3B", x"3B", x"37", x"32", x"00", x"00", x"00"),
(x"2E", x"37", x"3B", x"37", x"37", x"37", x"3B", x"3B", x"32", x"32", x"37", x"33", x"29", x"29", x"25", x"24", x"25", x"25", x"29", x"29", x"29", x"29", x"2E", x"32", x"37", x"32", x"2E", x"29", x"29", x"25", x"29", x"33", x"37", x"37", x"37", x"37", x"33", x"37", x"37", x"37", x"37", x"04", x"00", x"00"),
(x"2E", x"37", x"37", x"37", x"3B", x"37", x"37", x"33", x"2E", x"2D", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"3B", x"3B", x"32", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"32", x"2E", x"32", x"37", x"37", x"29", x"04", x"00"),
(x"32", x"37", x"37", x"3B", x"37", x"29", x"29", x"25", x"24", x"24", x"2E", x"37", x"3B", x"3B", x"3B", x"3B", x"3B", x"3B", x"3B", x"3B", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"32", x"37", x"37", x"37", x"33", x"33", x"32", x"37", x"37", x"37", x"2E", x"29"),
(x"32", x"3B", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"3B", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E"),
(x"32", x"3B", x"3B", x"37", x"25", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"3B", x"37", x"37", x"3B", x"37", x"37", x"37", x"37", x"37", x"32"),
(x"33", x"3B", x"3B", x"32", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"25", x"37", x"3B", x"37", x"37", x"37", x"37", x"37", x"3B", x"37", x"37", x"32"),
(x"33", x"3B", x"3B", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"25", x"33", x"3B", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"3B", x"33"),
(x"33", x"3B", x"3B", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"25", x"33", x"3B", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"3B", x"33"),
(x"33", x"3B", x"3B", x"32", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"25", x"37", x"3B", x"37", x"37", x"37", x"37", x"37", x"3B", x"37", x"37", x"32"),
(x"32", x"3B", x"3B", x"37", x"25", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"3B", x"37", x"37", x"3B", x"37", x"37", x"37", x"37", x"37", x"32"),
(x"32", x"3B", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"3B", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"2E"),
(x"32", x"37", x"37", x"3B", x"37", x"29", x"29", x"25", x"24", x"24", x"2E", x"37", x"3B", x"3B", x"3B", x"3B", x"3B", x"3B", x"3B", x"3B", x"37", x"37", x"37", x"37", x"2E", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"32", x"37", x"37", x"37", x"33", x"33", x"32", x"37", x"37", x"37", x"2E", x"29"),
(x"2E", x"37", x"37", x"37", x"3B", x"37", x"37", x"33", x"2E", x"2D", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"3B", x"3B", x"32", x"24", x"24", x"24", x"24", x"24", x"24", x"29", x"37", x"37", x"37", x"37", x"32", x"2E", x"32", x"37", x"37", x"29", x"04", x"00"),
(x"2E", x"37", x"3B", x"37", x"37", x"37", x"3B", x"3B", x"32", x"32", x"37", x"33", x"29", x"29", x"25", x"24", x"25", x"25", x"29", x"29", x"29", x"29", x"2E", x"32", x"37", x"32", x"2E", x"29", x"29", x"25", x"29", x"33", x"37", x"37", x"37", x"37", x"33", x"37", x"37", x"37", x"37", x"04", x"00", x"00"),
(x"29", x"33", x"37", x"37", x"3B", x"3B", x"3B", x"37", x"37", x"37", x"37", x"37", x"32", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"2E", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"3B", x"3B", x"37", x"32", x"00", x"00", x"00"),
(x"00", x"09", x"2D", x"2E", x"33", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"33", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"37", x"32", x"29", x"00", x"00", x"00"),
(x"00", x"00", x"20", x"00", x"04", x"09", x"29", x"2E", x"2E", x"2E", x"2E", x"2E", x"2E", x"2E", x"2D", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"29", x"09", x"33", x"32", x"05", x"29", x"29", x"29", x"29", x"2E", x"2E", x"2E", x"2E", x"2E", x"2E", x"29", x"00", x"2D", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"2E", x"29", x"37", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("00000000011000000000000011100000011110000000"),
("00011111111111111111111111111111111111110000"),
("11111111111111111111111111111111111111111100"),
("11111111111111111111111111111111111111111110"),
("11111111111111111111111111111111111111111110"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111110"),
("11111111111111111111111111111111111111111110"),
("11111111111111111111111111111111111111111100"),
("00011111111111111111111111111111111111110000"),
("00000000011000000000000011100000011110000000")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;
  end process;
end behav;		

--generated with PNGtoVHDL tool by Ben Wellingstein
