library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity restartEnter150X17_object is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end restartEnter150X17_object;

architecture behav of restartEnter150X17_object is

constant object_X_size : integer := 150;
constant object_Y_size : integer := 17;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"0C", x"76", x"DF", x"DF", x"DF", x"DF", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"9A", x"DF", x"DF", x"DF", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C"),
(x"0C", x"9A", x"FF", x"9A", x"96", x"96", x"DF", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"FF", x"96", x"96", x"96", x"51", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"55", x"FF", x"31", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"BA", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"31", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"11", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"11", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"31", x"0C", x"0C", x"0C", x"55", x"FF", x"31", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"BA", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"51", x"FF", x"31", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"BA", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"51", x"DF", x"31", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"BA", x"BB", x"0C", x"0C", x"0D", x"0C", x"0C", x"0D", x"0C", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"0C", x"0C", x"0D", x"0C", x"0C", x"0C", x"76", x"DF", x"31", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0D", x"0C", x"0C", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"BB", x"9A", x"0D", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"0C", x"0C", x"0D", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0D", x"BB", x"9A", x"0D", x"0C", x"0C", x"0C", x"0D", x"0D", x"0D", x"0D", x"0C", x"0C", x"0C", x"0D", x"0C", x"0C", x"0D", x"0C", x"0C", x"55", x"FF", x"31", x"0C", x"0C", x"51", x"DF", x"31", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"BA", x"BB", x"0C", x"0C", x"BA", x"BA", x"9A", x"DB", x"BA", x"0D", x"11", x"BA", x"DF", x"DF", x"DF", x"BB", x"31", x"0C", x"31", x"DB", x"DF", x"DF", x"DF", x"9A", x"0D", x"0C", x"76", x"DF", x"DF", x"DF", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"76", x"BB", x"96", x"BA", x"DB", x"BA", x"0C", x"51", x"DF", x"FF", x"DF", x"76", x"0C", x"55", x"DF", x"DF", x"DF", x"DF", x"96", x"0C", x"0D", x"BA", x"BA", x"BA", x"DB", x"9A", x"0C", x"0C", x"0C", x"0C", x"0C", x"9A", x"FF", x"FF", x"BB", x"31", x"0C", x"9A", x"DF", x"DF", x"DF", x"DB", x"51", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"DB", x"9A", x"BB", x"DF", x"55", x"0C", x"55", x"DF", x"DF", x"DF", x"DF", x"96", x"0C", x"0C", x"96", x"DF", x"DF", x"DF", x"DF", x"55", x"0C", x"9A", x"FF", x"FF", x"BB", x"31", x"0C", x"76", x"DF", x"DF", x"DF", x"DB", x"31", x"0C", x"51", x"DB", x"9A", x"BB", x"DF", x"51", x"51", x"DF", x"FF", x"DF", x"76", x"0C", x"51", x"DF", x"31", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"BA", x"BB", x"0C", x"0D", x"DB", x"DF", x"76", x"76", x"DF", x"11", x"31", x"FF", x"76", x"31", x"51", x"DF", x"51", x"0C", x"76", x"DF", x"51", x"31", x"76", x"DF", x"11", x"0C", x"BB", x"BA", x"31", x"31", x"9A", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"FF", x"9A", x"9A", x"9A", x"31", x"0C", x"76", x"FF", x"9A", x"76", x"76", x"DF", x"11", x"0D", x"96", x"FF", x"55", x"31", x"0C", x"9A", x"DB", x"51", x"31", x"96", x"DF", x"0D", x"0D", x"DF", x"DB", x"76", x"96", x"DF", x"0D", x"0C", x"0C", x"0C", x"0C", x"31", x"DF", x"BA", x"31", x"0C", x"31", x"DF", x"76", x"31", x"51", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"FF", x"9A", x"76", x"BB", x"9A", x"0C", x"9A", x"DB", x"51", x"31", x"96", x"DF", x"0D", x"0D", x"DF", x"9A", x"31", x"51", x"BB", x"9A", x"0C", x"31", x"DF", x"BA", x"31", x"0D", x"0C", x"DB", x"9A", x"31", x"51", x"DF", x"76", x"0C", x"55", x"FF", x"9A", x"76", x"DB", x"96", x"0D", x"76", x"FF", x"56", x"31", x"0C", x"31", x"DF", x"31", x"0C"),
(x"0C", x"9A", x"FF", x"9A", x"96", x"96", x"DF", x"BB", x"0C", x"0C", x"DB", x"76", x"0C", x"31", x"DF", x"11", x"31", x"FF", x"31", x"0C", x"0D", x"DF", x"55", x"0C", x"76", x"DF", x"0C", x"0C", x"31", x"DF", x"11", x"0C", x"BB", x"9A", x"0C", x"0C", x"76", x"BA", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"FF", x"BB", x"BB", x"BA", x"31", x"0C", x"76", x"DB", x"0C", x"0C", x"31", x"DF", x"11", x"0C", x"55", x"DF", x"0D", x"0C", x"0C", x"9A", x"BA", x"0C", x"0C", x"55", x"DF", x"0D", x"0D", x"DF", x"76", x"0C", x"51", x"DF", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"9A", x"9A", x"0C", x"9A", x"BA", x"0C", x"0C", x"55", x"DF", x"0D", x"0D", x"DF", x"76", x"0C", x"0C", x"9A", x"9A", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"0C", x"BA", x"76", x"0C", x"0C", x"BB", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"BA", x"96", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"31", x"DF", x"31", x"0C"),
(x"0C", x"9A", x"FF", x"DF", x"DB", x"DB", x"DB", x"76", x"0C", x"0D", x"DB", x"76", x"0C", x"31", x"76", x"0D", x"31", x"FF", x"31", x"0C", x"0D", x"DF", x"55", x"0C", x"51", x"FF", x"76", x"0C", x"0C", x"31", x"0C", x"0C", x"96", x"DF", x"51", x"0C", x"11", x"31", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"76", x"DB", x"0D", x"0C", x"31", x"DF", x"11", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"9A", x"BA", x"0C", x"0C", x"76", x"DF", x"0D", x"0D", x"DF", x"76", x"0C", x"31", x"76", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"55", x"55", x"0C", x"9A", x"BA", x"0C", x"0C", x"76", x"DF", x"0D", x"0C", x"BA", x"DF", x"31", x"0C", x"31", x"31", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"0C", x"0D", x"0D", x"0C", x"0D", x"BB", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"76", x"51", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"31", x"DF", x"11", x"0C"),
(x"0C", x"9A", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"DB", x"76", x"0C", x"0C", x"0C", x"0C", x"31", x"FF", x"DB", x"BB", x"BB", x"FF", x"51", x"0C", x"0C", x"56", x"DF", x"9A", x"11", x"0C", x"0C", x"0C", x"0D", x"96", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"76", x"DB", x"0D", x"0C", x"31", x"DF", x"11", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"9A", x"FF", x"BB", x"BB", x"DF", x"DB", x"0C", x"0D", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"0C", x"0C", x"9A", x"FF", x"BB", x"BB", x"DF", x"DB", x"0D", x"0C", x"11", x"BA", x"DF", x"56", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"0C", x"76", x"BB", x"BB", x"BB", x"FF", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"31", x"DB", x"11", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"DB", x"76", x"0C", x"0C", x"0C", x"0C", x"31", x"FF", x"76", x"55", x"56", x"55", x"0D", x"0C", x"0C", x"0C", x"31", x"DF", x"BB", x"31", x"0C", x"0C", x"0C", x"0C", x"76", x"DF", x"9A", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"76", x"DB", x"0D", x"0C", x"31", x"DF", x"11", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"9A", x"DF", x"76", x"56", x"56", x"31", x"0C", x"0D", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"0C", x"0C", x"9A", x"DF", x"76", x"56", x"56", x"31", x"0C", x"0C", x"0C", x"0C", x"76", x"FF", x"96", x"0D", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"9A", x"55", x"76", x"DF", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"31", x"BB", x"0D", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"DB", x"76", x"0C", x"0C", x"0C", x"0C", x"31", x"FF", x"31", x"0C", x"0C", x"0D", x"0C", x"0C", x"11", x"31", x"0C", x"31", x"BB", x"DB", x"0D", x"0C", x"31", x"11", x"0C", x"51", x"DF", x"9A", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"76", x"DB", x"0D", x"0C", x"31", x"DF", x"11", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"9A", x"BA", x"0C", x"0C", x"0C", x"0D", x"0C", x"0D", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"0C", x"0C", x"9A", x"BA", x"0C", x"0C", x"0C", x"0D", x"0C", x"0C", x"31", x"0D", x"0C", x"55", x"DF", x"76", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"11", x"76", x"0D", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"DB", x"76", x"0C", x"0C", x"0C", x"0C", x"31", x"FF", x"31", x"0C", x"0D", x"BA", x"51", x"0C", x"76", x"BB", x"0C", x"0C", x"51", x"DF", x"11", x"0C", x"BB", x"96", x"0C", x"0C", x"76", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"76", x"DB", x"0D", x"0C", x"31", x"DF", x"11", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"9A", x"BA", x"0C", x"0C", x"51", x"BA", x"0C", x"0D", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"0C", x"0C", x"9A", x"BA", x"0C", x"0C", x"51", x"BA", x"0C", x"0D", x"DB", x"76", x"0C", x"0C", x"9A", x"9A", x"0C", x"0C", x"BB", x"96", x"0C", x"0C", x"31", x"DF", x"51", x"0C", x"0C", x"BB", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C"),
(x"0C", x"9A", x"DF", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"DB", x"76", x"0C", x"0C", x"0C", x"0C", x"31", x"FF", x"51", x"0D", x"31", x"DF", x"55", x"0C", x"76", x"DF", x"31", x"0D", x"51", x"DF", x"11", x"0C", x"BB", x"9A", x"0D", x"0D", x"96", x"BB", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"DF", x"51", x"31", x"31", x"11", x"0C", x"76", x"DB", x"0D", x"0C", x"31", x"DF", x"11", x"0C", x"55", x"DF", x"31", x"0D", x"0C", x"9A", x"BB", x"11", x"0D", x"76", x"DF", x"0D", x"0D", x"DF", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"9A", x"0D", x"0C", x"31", x"DF", x"56", x"0D", x"31", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"0C", x"0C", x"9A", x"BB", x"11", x"0D", x"76", x"DF", x"0D", x"0D", x"DF", x"76", x"0D", x"11", x"BA", x"9A", x"0C", x"0C", x"BB", x"9A", x"0D", x"0C", x"31", x"DF", x"76", x"31", x"55", x"DF", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"51", x"FF", x"31", x"0D", x"0C", x"31", x"9A", x"31", x"0C"),
(x"0C", x"9A", x"DB", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BB", x"76", x"0C", x"0C", x"0C", x"0C", x"31", x"DF", x"DF", x"DF", x"DF", x"DF", x"31", x"0C", x"51", x"DF", x"DF", x"DF", x"DF", x"BB", x"0D", x"0C", x"96", x"DF", x"DF", x"DF", x"DF", x"96", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"BA", x"FF", x"FF", x"FF", x"FF", x"76", x"0C", x"76", x"BB", x"0C", x"0C", x"31", x"DF", x"11", x"0C", x"31", x"DF", x"DF", x"76", x"0C", x"76", x"DF", x"DF", x"DF", x"DF", x"BA", x"0C", x"0D", x"DB", x"76", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"96", x"DF", x"DB", x"31", x"0D", x"BB", x"DF", x"DF", x"DF", x"DF", x"55", x"0C", x"0C", x"0C", x"0C", x"0C", x"51", x"DF", x"31", x"0C", x"0C", x"0C", x"0C", x"76", x"DF", x"DF", x"DF", x"DF", x"BA", x"0C", x"0C", x"9A", x"DF", x"DF", x"DF", x"DF", x"76", x"0C", x"0C", x"96", x"DF", x"DB", x"31", x"0D", x"BB", x"DF", x"DF", x"BB", x"DF", x"76", x"0C", x"55", x"DF", x"11", x"0C", x"0C", x"0C", x"0C", x"31", x"DF", x"DF", x"76", x"0C", x"55", x"FF", x"31", x"0C"),
(x"0C", x"31", x"31", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"11", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"31", x"31", x"31", x"31", x"0C", x"0C", x"0C", x"31", x"31", x"31", x"31", x"11", x"0C", x"0C", x"0D", x"31", x"31", x"31", x"31", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"31", x"31", x"31", x"31", x"11", x"0C", x"11", x"31", x"0C", x"0C", x"0D", x"31", x"0C", x"0C", x"0C", x"31", x"31", x"31", x"0C", x"0C", x"31", x"31", x"31", x"31", x"11", x"0C", x"0C", x"31", x"0D", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"31", x"31", x"0D", x"0C", x"11", x"31", x"31", x"31", x"31", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"0D", x"31", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"31", x"31", x"31", x"11", x"0C", x"0C", x"0D", x"31", x"31", x"31", x"31", x"0D", x"0C", x"0C", x"0D", x"31", x"31", x"0D", x"0C", x"31", x"31", x"31", x"0D", x"31", x"11", x"0C", x"0D", x"31", x"0C", x"0C", x"0C", x"0C", x"0C", x"0C", x"31", x"31", x"31", x"0C", x"0D", x"31", x"0D", x"0C")
);

-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;
  end process;
end behav;		

--generated with PNGtoVHDL tool by Ben Wellingstein
