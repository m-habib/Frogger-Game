library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity plank_141_30_object is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end plank_141_30_object;

architecture behav of plank_141_30_object is

constant object_X_size : integer := 141;
constant object_Y_size : integer := 30;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"20", x"64", x"64", x"64", x"64", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"88", x"88", x"64", x"64", x"44", x"44", x"44", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"88", x"88", x"68", x"91", x"B1", x"6D", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"D5", x"FA", x"FA", x"FA", x"69", x"00", x"00"),
(x"00", x"00", x"00", x"20", x"88", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"AD", x"FA", x"FA", x"F6", x"F6", x"B1", x"20", x"00"),
(x"00", x"00", x"00", x"64", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"A8", x"D1", x"FA", x"FA", x"FA", x"FA", x"F6", x"48", x"00"),
(x"00", x"00", x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"D6", x"F6", x"FA", x"F6", x"FA", x"F6", x"69", x"00"),
(x"00", x"00", x"64", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"8C", x"F6", x"F6", x"FA", x"FA", x"F6", x"F6", x"8D", x"00"),
(x"00", x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"8D", x"FA", x"F6", x"FA", x"FA", x"FA", x"FA", x"8D", x"00"),
(x"00", x"44", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"B1", x"FA", x"FA", x"FA", x"F6", x"F6", x"FA", x"B1", x"00"),
(x"00", x"64", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"B1", x"FA", x"FA", x"FA", x"F6", x"F6", x"FA", x"B1", x"00"),
(x"00", x"88", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"D1", x"FA", x"FA", x"FA", x"F6", x"F6", x"FA", x"B1", x"20"),
(x"20", x"A8", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"AC", x"D1", x"FA", x"FA", x"FA", x"F5", x"F6", x"F6", x"D1", x"20"),
(x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"D1", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"D1", x"20"),
(x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"B1", x"FA", x"FA", x"FA", x"F6", x"F5", x"F6", x"B1", x"20"),
(x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"AD", x"FA", x"FA", x"F6", x"F6", x"F5", x"F6", x"B1", x"00"),
(x"44", x"A8", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"AC", x"FA", x"FA", x"F6", x"F6", x"F6", x"FA", x"B1", x"00"),
(x"44", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"AC", x"D6", x"FA", x"F6", x"F6", x"F6", x"FA", x"B1", x"00"),
(x"44", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"AC", x"D5", x"FA", x"F6", x"F6", x"F6", x"F6", x"B1", x"00"),
(x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"B1", x"FA", x"F6", x"F6", x"FA", x"F6", x"B1", x"00"),
(x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"B1", x"FA", x"F6", x"F6", x"FA", x"FA", x"B1", x"00"),
(x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"AC", x"FA", x"F6", x"F6", x"F6", x"FA", x"D1", x"24"),
(x"00", x"88", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"AC", x"F6", x"FA", x"F6", x"F6", x"FA", x"D1", x"24"),
(x"00", x"64", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"AC", x"D6", x"F6", x"FA", x"F6", x"FA", x"B1", x"20"),
(x"00", x"44", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"D1", x"F6", x"FA", x"FA", x"FA", x"B1", x"00"),
(x"00", x"20", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"B1", x"FA", x"F6", x"FA", x"FA", x"8D", x"00"),
(x"00", x"00", x"88", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"AD", x"FA", x"F6", x"FA", x"FA", x"69", x"00"),
(x"00", x"00", x"64", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"C8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"8C", x"F6", x"FA", x"FA", x"D6", x"24", x"00"),
(x"00", x"00", x"20", x"88", x"A8", x"A8", x"88", x"64", x"64", x"44", x"44", x"44", x"64", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"A8", x"A8", x"A8", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"CC", x"A8", x"8D", x"D6", x"D6", x"68", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"44", x"44", x"44", x"44", x"20", x"20", x"20", x"20", x"20", x"20", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"64", x"64", x"64", x"64", x"64", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"20", x"24", x"24", x"00", x"00", x"00"),
(x"00", x"00", x"64", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"88", x"FC", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;
  end process;
end behav;		

--generated with PNGtoVHDL tool by Ben Wellingstein
