--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity WinsTable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(13 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end WinsTable;

architecture arch of WinsTable is
constant array_size 			: integer := 13926 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal Wins_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  WinsJumpTable_proc: process(resetN, CLK)
    constant Wins_table : table_type := (
---start 0 v

X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"0465",
X"03E8",
X"02EE",
X"0271",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"0465",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"07D0",
X"084D",
X"0947",
X"09C4",
X"0A41",
X"0ABE",
X"0BB8",
X"0C35",
X"0CB2",
X"0D2F",
X"0C35",
X"0BB8",
X"0B3B",
X"0ABE",
X"09C4",
X"0947",
X"084D",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"036B",
X"0465",
X"055F",
X"0659",
X"0753",
X"084D",
X"0947",
X"09C4",
X"0947",
X"08CA",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"06D6",
X"0659",
X"05DC",
X"04E2",
X"03E8",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F63C",
X"F5BF",
X"F5BF",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F542",
X"F5BF",
X"F63C",
X"F63C",
X"F6B9",
X"F736",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"06D6",
X"07D0",
X"084D",
X"08CA",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"0465",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F7B3",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"0465",
X"055F",
X"0659",
X"0753",
X"084D",
X"0947",
X"09C4",
X"0947",
X"08CA",
X"08CA",
X"084D",
X"07D0",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0BB8",
X"0C35",
X"0CB2",
X"0C35",
X"0B3B",
X"0A41",
X"0947",
X"084D",
X"0753",
X"0659",
X"055F",
X"0465",
X"036B",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"06D6",
X"0753",
X"084D",
X"08CA",
X"0947",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0C35",
X"0CB2",
X"0C35",
X"0B3B",
X"0ABE",
X"0A41",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F7B3",
X"F736",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"0659",
X"0753",
X"084D",
X"0947",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0BB8",
X"0C35",
X"0CB2",
X"0BB8",
X"0ABE",
X"0947",
X"084D",
X"0753",
X"0659",
X"055F",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"0659",
X"0753",
X"084D",
X"08CA",
X"09C4",
X"0A41",
X"0ABE",
X"0BB8",
X"0C35",
X"0CB2",
X"0CB2",
X"0C35",
X"0B3B",
X"0ABE",
X"09C4",
X"0947",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"05DC",
X"06D6",
X"084D",
X"0947",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"06D6",
X"0659",
X"055F",
X"03E8",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F63C",
X"F5BF",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F5BF",
X"F63C",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"036B",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"0753",
X"07D0",
X"08CA",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"0659",
X"07D0",
X"08CA",
X"09C4",
X"0947",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"09C4",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0C35",
X"0C35",
X"0C35",
X"0B3B",
X"0A41",
X"0947",
X"084D",
X"06D6",
X"05DC",
X"04E2",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F7B3",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"02EE",
X"03E8",
X"04E2",
X"0659",
X"0753",
X"08CA",
X"09C4",
X"0947",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0BB8",
X"0C35",
X"0CB2",
X"0B3B",
X"0A41",
X"0947",
X"07D0",
X"06D6",
X"05DC",
X"0465",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"0659",
X"0753",
X"084D",
X"08CA",
X"09C4",
X"0A41",
X"0B3B",
X"0BB8",
X"0CB2",
X"0D2F",
X"0C35",
X"0BB8",
X"0ABE",
X"0A41",
X"0947",
X"084D",
X"07D0",
X"06D6",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"0177",
X"0271",
X"036B",
X"0465",
X"05DC",
X"06D6",
X"07D0",
X"08CA",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"055F",
X"0465",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FE89",
X"FD8F",
X"FC95",
X"FC18",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F542",
X"F5BF",
X"F63C",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0271",
X"036B",
X"03E8",
X"04E2",
X"05DC",
X"0659",
X"0753",
X"07D0",
X"08CA",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"036B",
X"0465",
X"05DC",
X"06D6",
X"07D0",
X"0947",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"0177",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0C35",
X"0CB2",
X"0C35",
X"0ABE",
X"09C4",
X"08CA",
X"0753",
X"0659",
X"055F",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"0753",
X"07D0",
X"084D",
X"0947",
X"09C4",
X"0A41",
X"0ABE",
X"0B3B",
X"0B3B",
X"0A41",
X"09C4",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"02EE",
X"03E8",
X"04E2",
X"0659",
X"0753",
X"08CA",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"05DC",
X"0465",
X"036B",
X"01F4",
X"007D",
X"FF83",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"05DC",
X"06D6",
X"0753",
X"084D",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"04E2",
X"0465",
X"036B",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"036B",
X"04E2",
X"0659",
X"0753",
X"08CA",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0ABE",
X"0B3B",
X"0BB8",
X"0C35",
X"0CB2",
X"0C35",
X"0ABE",
X"09C4",
X"084D",
X"06D6",
X"05DC",
X"0465",
X"036B",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"06D6",
X"07D0",
X"08CA",
X"09C4",
X"0A41",
X"0B3B",
X"0C35",
X"0CB2",
X"0CB2",
X"0BB8",
X"0B3B",
X"0A41",
X"0947",
X"084D",
X"0753",
X"0659",
X"055F",
X"055F",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"00FA",
X"01F4",
X"036B",
X"0465",
X"05DC",
X"06D6",
X"084D",
X"0947",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"05DC",
X"0465",
X"036B",
X"01F4",
X"007D",
X"FF83",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"05DC",
X"06D6",
X"0753",
X"084D",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"036B",
X"04E2",
X"0659",
X"0753",
X"08CA",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"0465",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0659",
X"04E2",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F63C",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"0659",
X"0753",
X"084D",
X"08CA",
X"084D",
X"0753",
X"0659",
X"05DC",
X"04E2",
X"036B",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"0000",
X"0177",
X"02EE",
X"0465",
X"05DC",
X"0753",
X"08CA",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"036B",
X"03E8",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0B3B",
X"0BB8",
X"0C35",
X"0CB2",
X"0BB8",
X"0A41",
X"08CA",
X"0753",
X"05DC",
X"0465",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"06D6",
X"07D0",
X"08CA",
X"09C4",
X"0ABE",
X"0BB8",
X"0C35",
X"0D2F",
X"0C35",
X"0B3B",
X"0A41",
X"0947",
X"084D",
X"0753",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"036B",
X"02EE",
X"0271",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"00FA",
X"01F4",
X"036B",
X"04E2",
X"0659",
X"07D0",
X"0947",
X"09C4",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"055F",
X"03E8",
X"0271",
X"00FA",
X"FF83",
X"FE0C",
X"FD12",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F736",
X"F6B9",
X"F63C",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0271",
X"036B",
X"04E2",
X"05DC",
X"06D6",
X"07D0",
X"08CA",
X"08CA",
X"07D0",
X"06D6",
X"05DC",
X"055F",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FAA1",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"036B",
X"04E2",
X"0659",
X"07D0",
X"0947",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"09C4",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0C35",
X"0C35",
X"0ABE",
X"0947",
X"07D0",
X"0659",
X"04E2",
X"036B",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"0753",
X"084D",
X"0947",
X"0A41",
X"0B3B",
X"0C35",
X"0CB2",
X"0CB2",
X"0BB8",
X"0ABE",
X"09C4",
X"08CA",
X"07D0",
X"0659",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"0659",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"04E2",
X"05DC",
X"0659",
X"0753",
X"07D0",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"04E2",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"0271",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0177",
X"02EE",
X"0465",
X"05DC",
X"0753",
X"0947",
X"09C4",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FC95",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"055F",
X"03E8",
X"0271",
X"007D",
X"FF06",
X"FD8F",
X"FC18",
X"FB9B",
X"FAA1",
X"F9A7",
X"F92A",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F92A",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"036B",
X"0465",
X"055F",
X"06D6",
X"07D0",
X"08CA",
X"084D",
X"0753",
X"0659",
X"055F",
X"0465",
X"036B",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F92A",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"055F",
X"0753",
X"08CA",
X"09C4",
X"0947",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"0A41",
X"0ABE",
X"0B3B",
X"0C35",
X"0CB2",
X"0B3B",
X"09C4",
X"084D",
X"0659",
X"04E2",
X"036B",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"0753",
X"08CA",
X"09C4",
X"0ABE",
X"0BB8",
X"0CB2",
X"0CB2",
X"0BB8",
X"0ABE",
X"0947",
X"084D",
X"06D6",
X"05DC",
X"055F",
X"0465",
X"03E8",
X"036B",
X"0271",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"055F",
X"06D6",
X"08CA",
X"09C4",
X"0947",
X"084D",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"0659",
X"06D6",
X"05DC",
X"0465",
X"0271",
X"00FA",
X"FF83",
X"FE0C",
X"FC95",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F8AD",
X"F7B3",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F542",
X"F5BF",
X"F63C",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"0177",
X"02EE",
X"03E8",
X"055F",
X"0659",
X"0753",
X"084D",
X"08CA",
X"07D0",
X"06D6",
X"05DC",
X"0465",
X"036B",
X"0271",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"01F4",
X"036B",
X"04E2",
X"06D6",
X"084D",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0ABE",
X"0B3B",
X"0BB8",
X"0CB2",
X"0BB8",
X"0A41",
X"08CA",
X"06D6",
X"055F",
X"03E8",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0753",
X"084D",
X"0947",
X"0A41",
X"0B3B",
X"0C35",
X"0CB2",
X"0BB8",
X"0ABE",
X"09C4",
X"084D",
X"0753",
X"0659",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"0465",
X"05DC",
X"06D6",
X"084D",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"007D",
X"0177",
X"02EE",
X"0465",
X"05DC",
X"0753",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"03E8",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"0A41",
X"0ABE",
X"0B3B",
X"0C35",
X"0CB2",
X"0B3B",
X"0947",
X"07D0",
X"05DC",
X"0465",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0753",
X"084D",
X"09C4",
X"0ABE",
X"0BB8",
X"0CB2",
X"0CB2",
X"0B3B",
X"0A41",
X"08CA",
X"07D0",
X"0659",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"036B",
X"055F",
X"06D6",
X"08CA",
X"09C4",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FC95",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"04E2",
X"055F",
X"05DC",
X"06D6",
X"05DC",
X"0465",
X"0271",
X"00FA",
X"FF06",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F8AD",
X"F830",
X"F7B3",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"0177",
X"0271",
X"036B",
X"04E2",
X"05DC",
X"0753",
X"084D",
X"08CA",
X"07D0",
X"06D6",
X"05DC",
X"0465",
X"036B",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"00FA",
X"0271",
X"0465",
X"0659",
X"07D0",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"0465",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"09C4",
X"0A41",
X"0ABE",
X"0BB8",
X"0C35",
X"0C35",
X"0ABE",
X"08CA",
X"0753",
X"055F",
X"03E8",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"0177",
X"0271",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"0659",
X"0753",
X"08CA",
X"09C4",
X"0ABE",
X"0BB8",
X"0D2F",
X"0C35",
X"0B3B",
X"09C4",
X"08CA",
X"0753",
X"0659",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0271",
X"03E8",
X"05DC",
X"0753",
X"08CA",
X"09C4",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FC95",
X"FB9B",
X"FAA1",
X"F9A7",
X"F92A",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"0659",
X"06D6",
X"05DC",
X"03E8",
X"01F4",
X"007D",
X"FF06",
X"FD12",
X"FC18",
X"FB1E",
X"FA24",
X"F9A7",
X"F8AD",
X"F830",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F92A",
X"F9A7",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"03E8",
X"04E2",
X"0659",
X"0753",
X"084D",
X"08CA",
X"07D0",
X"0659",
X"055F",
X"0465",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F7B3",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"0177",
X"02EE",
X"04E2",
X"0659",
X"084D",
X"09C4",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"06D6",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"0465",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"09C4",
X"0A41",
X"0B3B",
X"0BB8",
X"0C35",
X"0C35",
X"0A41",
X"08CA",
X"06D6",
X"055F",
X"036B",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"07D0",
X"08CA",
X"0A41",
X"0B3B",
X"0C35",
X"0D2F",
X"0C35",
X"0ABE",
X"09C4",
X"084D",
X"0753",
X"05DC",
X"055F",
X"0465",
X"03E8",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"02EE",
X"0465",
X"05DC",
X"07D0",
X"0947",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD12",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"06D6",
X"055F",
X"036B",
X"01F4",
X"0000",
X"FE89",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F92A",
X"F8AD",
X"F7B3",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F92A",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"02EE",
X"03E8",
X"055F",
X"0659",
X"07D0",
X"08CA",
X"084D",
X"0753",
X"0659",
X"055F",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F92A",
X"F9A7",
X"FA24",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"0000",
X"0177",
X"036B",
X"04E2",
X"06D6",
X"08CA",
X"09C4",
X"0947",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0ABE",
X"0B3B",
X"0BB8",
X"0CB2",
X"0BB8",
X"09C4",
X"084D",
X"0659",
X"04E2",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"06D6",
X"07D0",
X"0947",
X"0A41",
X"0B3B",
X"0C35",
X"0CB2",
X"0BB8",
X"0ABE",
X"0947",
X"084D",
X"06D6",
X"05DC",
X"04E2",
X"0465",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"0177",
X"02EE",
X"04E2",
X"0659",
X"07D0",
X"09C4",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FD12",
X"FC18",
X"FB1E",
X"FA24",
X"F9A7",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"04E2",
X"02EE",
X"0177",
X"0000",
X"FE0C",
X"FC95",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F5BF",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"FA24",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"06D6",
X"07D0",
X"08CA",
X"084D",
X"0753",
X"05DC",
X"04E2",
X"03E8",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FAA1",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FE0C",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"055F",
X"0753",
X"08CA",
X"09C4",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0ABE",
X"0B3B",
X"0C35",
X"0CB2",
X"0B3B",
X"09C4",
X"07D0",
X"0659",
X"0465",
X"02EE",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"04E2",
X"055F",
X"05DC",
X"06D6",
X"084D",
X"0947",
X"0ABE",
X"0BB8",
X"0CB2",
X"0CB2",
X"0BB8",
X"0A41",
X"0947",
X"07D0",
X"06D6",
X"055F",
X"04E2",
X"0465",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"01F4",
X"036B",
X"04E2",
X"06D6",
X"084D",
X"09C4",
X"0947",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FD12",
X"FC18",
X"FB1E",
X"FA24",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"04E2",
X"055F",
X"05DC",
X"06D6",
X"0659",
X"0465",
X"02EE",
X"00FA",
X"FF83",
X"FD8F",
X"FC18",
X"FB9B",
X"FAA1",
X"F9A7",
X"F92A",
X"F830",
X"F7B3",
X"F736",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"0177",
X"01F4",
X"036B",
X"04E2",
X"05DC",
X"06D6",
X"084D",
X"08CA",
X"07D0",
X"06D6",
X"05DC",
X"04E2",
X"036B",
X"0271",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FC95",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FE0C",
X"FF06",
X"007D",
X"0271",
X"03E8",
X"05DC",
X"07D0",
X"0947",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"0659",
X"06D6",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"0A41",
X"0ABE",
X"0BB8",
X"0C35",
X"0CB2",
X"0ABE",
X"0947",
X"0753",
X"05DC",
X"03E8",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"007D",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0753",
X"084D",
X"09C4",
X"0ABE",
X"0BB8",
X"0CB2",
X"0C35",
X"0B3B",
X"0A41",
X"08CA",
X"07D0",
X"0659",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"055F",
X"0753",
X"08CA",
X"09C4",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FC95",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"0659",
X"06D6",
X"05DC",
X"03E8",
X"0271",
X"007D",
X"FF06",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F8AD",
X"F830",
X"F7B3",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F9A7",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"03E8",
X"04E2",
X"05DC",
X"0753",
X"084D",
X"08CA",
X"07D0",
X"06D6",
X"055F",
X"0465",
X"036B",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FE0C",
X"FF83",
X"00FA",
X"02EE",
X"0465",
X"0659",
X"07D0",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"0271",
X"036B",
X"0465",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"09C4",
X"0A41",
X"0ABE",
X"0BB8",
X"0C35",
X"0C35",
X"0ABE",
X"08CA",
X"0753",
X"055F",
X"03E8",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"0753",
X"08CA",
X"09C4",
X"0ABE",
X"0C35",
X"0D2F",
X"0C35",
X"0B3B",
X"09C4",
X"08CA",
X"0753",
X"0659",
X"055F",
X"0465",
X"03E8",
X"036B",
X"0271",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"05DC",
X"0753",
X"0947",
X"0947",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FC95",
X"FB9B",
X"FAA1",
X"F9A7",
X"F92A",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FB1E",
X"FC18",
X"FD12",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"06D6",
X"055F",
X"03E8",
X"01F4",
X"007D",
X"FE89",
X"FD12",
X"FC18",
X"FB1E",
X"FA24",
X"F9A7",
X"F8AD",
X"F830",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F92A",
X"F9A7",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"03E8",
X"055F",
X"0659",
X"0753",
X"08CA",
X"08CA",
X"0753",
X"0659",
X"055F",
X"0465",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F830",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FE89",
X"FF83",
X"0177",
X"02EE",
X"04E2",
X"06D6",
X"084D",
X"09C4",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"06D6",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"0465",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0B3B",
X"0BB8",
X"0C35",
X"0BB8",
X"0A41",
X"084D",
X"06D6",
X"04E2",
X"036B",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"0659",
X"07D0",
X"08CA",
X"0A41",
X"0B3B",
X"0C35",
X"0D2F",
X"0BB8",
X"0ABE",
X"09C4",
X"084D",
X"0753",
X"05DC",
X"055F",
X"0465",
X"03E8",
X"02EE",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"02EE",
X"0465",
X"0659",
X"07D0",
X"0947",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD12",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FE0C",
X"FF06",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"04E2",
X"036B",
X"0177",
X"0000",
X"FE89",
X"FC95",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F8AD",
X"F7B3",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F6B9",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F92A",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"0177",
X"02EE",
X"0465",
X"055F",
X"06D6",
X"07D0",
X"08CA",
X"084D",
X"0753",
X"0659",
X"04E2",
X"03E8",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"0000",
X"01F4",
X"036B",
X"055F",
X"06D6",
X"08CA",
X"09C4",
X"0947",
X"084D",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"0271",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0ABE",
X"0B3B",
X"0BB8",
X"0CB2",
X"0BB8",
X"09C4",
X"084D",
X"0659",
X"04E2",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"04E2",
X"055F",
X"05DC",
X"06D6",
X"07D0",
X"0947",
X"0A41",
X"0B3B",
X"0CB2",
X"0CB2",
X"0BB8",
X"0ABE",
X"0947",
X"084D",
X"06D6",
X"05DC",
X"04E2",
X"0465",
X"036B",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"0177",
X"036B",
X"04E2",
X"0659",
X"084D",
X"09C4",
X"0947",
X"084D",
X"07D0",
X"0753",
X"0659",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD12",
X"FD12",
X"FC18",
X"FB1E",
X"FA24",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB9B",
X"FC95",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"0659",
X"0659",
X"04E2",
X"02EE",
X"0177",
X"FF83",
X"FE0C",
X"FC95",
X"FB9B",
X"FAA1",
X"F9A7",
X"F92A",
X"F830",
X"F7B3",
X"F736",
X"F63C",
X"F5BF",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F63C",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F9A7",
X"FA24",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"036B",
X"0465",
X"05DC",
X"06D6",
X"07D0",
X"08CA",
X"084D",
X"06D6",
X"05DC",
X"04E2",
X"036B",
X"0271",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FAA1",
X"FB9B",
X"FC18",
X"FD12",
X"FE0C",
X"FF06",
X"007D",
X"01F4",
X"03E8",
X"055F",
X"0753",
X"0947",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"00FA",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"0947",
X"09C4",
X"0A41",
X"0B3B",
X"0BB8",
X"0C35",
X"0ABE",
X"0947",
X"0753",
X"05DC",
X"0465",
X"0271",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"0465",
X"055F",
X"05DC",
X"06D6",
X"07D0",
X"0947",
X"0A41",
X"0B3B",
X"0C35",
X"0C35",
X"0ABE",
X"09C4",
X"08CA",
X"0753",
X"0659",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"007D",
X"01F4",
X"036B",
X"04E2",
X"0659",
X"07D0",
X"0947",
X"084D",
X"07D0",
X"0753",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FD12",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC18",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"0659",
X"055F",
X"03E8",
X"0271",
X"00FA",
X"FF83",
X"FD8F",
X"FC95",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F5BF",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"FA24",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"0659",
X"0753",
X"07D0",
X"0753",
X"0659",
X"055F",
X"03E8",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F8AD",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FF06",
X"007D",
X"0271",
X"03E8",
X"055F",
X"06D6",
X"084D",
X"084D",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF83",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"0753",
X"0753",
X"07D0",
X"084D",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0ABE",
X"0947",
X"07D0",
X"0659",
X"04E2",
X"036B",
X"01F4",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"0659",
X"0753",
X"084D",
X"0947",
X"0A41",
X"0ABE",
X"0A41",
X"0947",
X"084D",
X"0753",
X"0659",
X"055F",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE0C",
X"FE89",
X"FF83",
X"007D",
X"01F4",
X"036B",
X"0465",
X"05DC",
X"0753",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"04E2",
X"0465",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC95",
X"FD12",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC95",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"0465",
X"036B",
X"01F4",
X"007D",
X"FF06",
X"FD8F",
X"FC95",
X"FC18",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"05DC",
X"06D6",
X"06D6",
X"05DC",
X"055F",
X"0465",
X"036B",
X"0271",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"00FA",
X"0271",
X"036B",
X"04E2",
X"0659",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"06D6",
X"0753",
X"07D0",
X"084D",
X"08CA",
X"0947",
X"0947",
X"07D0",
X"0659",
X"055F",
X"03E8",
X"0271",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"0753",
X"084D",
X"08CA",
X"09C4",
X"08CA",
X"084D",
X"0753",
X"0659",
X"055F",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"01F4",
X"02EE",
X"0465",
X"055F",
X"06D6",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"03E8",
X"0271",
X"0177",
X"0000",
X"FF06",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"0465",
X"055F",
X"05DC",
X"05DC",
X"04E2",
X"0465",
X"036B",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"036B",
X"0465",
X"05DC",
X"0659",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"007D",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"0659",
X"06D6",
X"0753",
X"07D0",
X"084D",
X"07D0",
X"0659",
X"055F",
X"0465",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"036B",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"0753",
X"07D0",
X"084D",
X"0753",
X"06D6",
X"05DC",
X"055F",
X"0465",
X"036B",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"05DC",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"03E8",
X"02EE",
X"01F4",
X"00FA",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0271",
X"02EE",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"06D6",
X"0659",
X"055F",
X"0465",
X"036B",
X"0271",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"06D6",
X"06D6",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"0271",
X"036B",
X"0465",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"036B",
X"03E8",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"01F4",
X"0271",
X"036B",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"0271",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000"



 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= Wins_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;