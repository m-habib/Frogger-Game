library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity wood_object is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end wood_object;

architecture behav of wood_object is

constant object_X_size : integer := 115;
constant object_Y_size : integer := 30;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"44", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8D", x"91", x"88", x"8D", x"AD", x"AD", x"F6", x"D1", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8D", x"8D", x"8D", x"8D", x"89", x"8D", x"8D", x"8D", x"88", x"8D", x"8D", x"8D", x"B1", x"B2", x"92", x"91", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"AD", x"44", x"68", x"68", x"68", x"88", x"88", x"AC", x"AD", x"AD", x"AD", x"B1", x"D1", x"D1", x"D6", x"FF", x"FA", x"D1", x"AC", x"FF", x"D1", x"B1", x"AD", x"AD", x"8D", x"8C", x"88", x"8C", x"8C", x"8D", x"AD", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"AD", x"AD", x"B1", x"D6", x"B1", x"B1", x"B1", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"8D", x"8D", x"8D", x"8D", x"B6", x"FF", x"FF", x"00", x"00", x"00", x"00", x"D6", x"DA", x"FB", x"FB", x"FF", x"FF", x"B1", x"92", x"8D", x"FF", x"FF", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"D6", x"D6", x"D1", x"FA", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D1", x"00", x"88", x"64", x"44", x"64", x"88", x"AC", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"88", x"88", x"88", x"88", x"68", x"88", x"8D", x"AD", x"8D", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"89", x"8D", x"89", x"89", x"8D", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"89", x"8D", x"8D", x"8D", x"AD", x"AD", x"AD", x"8D", x"8D", x"8D", x"88", x"68", x"88", x"8D", x"AD", x"8D", x"8D", x"FF", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"FB", x"64", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8D", x"AD", x"AC", x"AC", x"AC", x"AC", x"AC", x"AD", x"AD", x"AC", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"AD", x"8C", x"8D", x"88", x"68", x"68", x"44", x"44", x"68", x"88", x"AC", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"8C", x"8C", x"8C", x"88", x"68", x"68", x"88", x"8C", x"88", x"8D", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8C", x"88", x"88", x"8D", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"88", x"89", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"89", x"88", x"88", x"88", x"68", x"88", x"89", x"89", x"8D", x"68", x"FF", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"D6", x"00", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8C", x"88", x"88", x"88", x"68", x"68", x"68", x"64", x"64", x"64", x"68", x"88", x"88", x"8C", x"8D", x"AD", x"8D", x"8D", x"8C", x"8C", x"8C", x"8C", x"8D", x"AD", x"8D", x"8C", x"8C", x"88", x"88", x"88", x"8C", x"88", x"88", x"68", x"44", x"44", x"88", x"88", x"88", x"88", x"8D", x"8D", x"AD", x"AD", x"8D", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"AD", x"AD", x"AD", x"AD", x"88", x"88", x"89", x"89", x"89", x"8D", x"8D", x"8D", x"8D", x"AD", x"AD", x"AD", x"8D", x"88", x"88", x"89", x"8D", x"8D", x"88", x"88", x"88", x"68", x"64", x"69", x"68", x"FF", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"8D", x"8D", x"68", x"68", x"88", x"68", x"68", x"68", x"88", x"88", x"68", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"64", x"64", x"64", x"68", x"68", x"68", x"88", x"88", x"88", x"68", x"64", x"44", x"44", x"68", x"88", x"88", x"88", x"AD", x"AD", x"AD", x"8D", x"8D", x"8C", x"8C", x"8C", x"8C", x"8C", x"8D", x"8D", x"8C", x"88", x"88", x"8C", x"8C", x"8C", x"8C", x"88", x"88", x"68", x"68", x"88", x"8D", x"8C", x"88", x"8C", x"8D", x"8D", x"8D", x"89", x"8D", x"8D", x"8D", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"AD", x"AD", x"8D", x"AD", x"AD", x"AD", x"8D", x"8D", x"88", x"8D", x"89", x"89", x"88", x"68", x"64", x"64", x"68", x"68", x"69", x"69", x"FF", x"00"),
(x"00", x"00", x"00", x"00", x"88", x"00", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"88", x"88", x"88", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"20", x"44", x"64", x"88", x"AD", x"AD", x"8D", x"8D", x"8D", x"8C", x"88", x"88", x"88", x"88", x"8C", x"AD", x"AD", x"8C", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"89", x"88", x"88", x"68", x"89", x"8D", x"88", x"64", x"68", x"68", x"68", x"69", x"68", x"FF", x"00"),
(x"00", x"00", x"00", x"FF", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"44", x"44", x"44", x"64", x"88", x"AD", x"AD", x"8D", x"8D", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8C", x"8C", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"AD", x"AD", x"AD", x"AD", x"8D", x"8D", x"8D", x"8D", x"88", x"88", x"8D", x"68", x"68", x"68", x"44", x"44", x"44", x"6D", x"69", x"FF", x"00"),
(x"00", x"00", x"00", x"FF", x"44", x"68", x"64", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"68", x"88", x"88", x"8C", x"8D", x"8C", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"8C", x"AD", x"88", x"88", x"68", x"68", x"68", x"68", x"88", x"8D", x"8D", x"8D", x"8D", x"88", x"88", x"88", x"88", x"8D", x"8D", x"8D", x"8D", x"8D", x"AD", x"AD", x"AD", x"8D", x"8D", x"89", x"89", x"89", x"89", x"89", x"89", x"89", x"88", x"68", x"64", x"44", x"44", x"20", x"20", x"44", x"44", x"44", x"48", x"20", x"6D", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"44", x"68", x"64", x"68", x"68", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"88", x"8C", x"8C", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"88", x"8C", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"68", x"88", x"88", x"88", x"68", x"88", x"88", x"88", x"8C", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"88", x"88", x"88", x"68", x"68", x"68", x"88", x"8D", x"8D", x"8D", x"89", x"89", x"8D", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"48", x"91", x"6D", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"44", x"44", x"44", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"8C", x"AD", x"AC", x"88", x"88", x"88", x"68", x"64", x"64", x"64", x"64", x"68", x"88", x"88", x"88", x"88", x"68", x"68", x"64", x"64", x"44", x"44", x"64", x"64", x"68", x"88", x"88", x"88", x"88", x"68", x"88", x"88", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"88", x"8C", x"88", x"68", x"68", x"88", x"89", x"89", x"8D", x"8D", x"8D", x"AD", x"AD", x"8D", x"88", x"68", x"68", x"64", x"44", x"44", x"68", x"00", x"B6", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"64", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8C", x"88", x"88", x"88", x"88", x"68", x"68", x"64", x"68", x"68", x"68", x"88", x"88", x"8C", x"88", x"88", x"88", x"68", x"68", x"64", x"64", x"64", x"68", x"68", x"88", x"8C", x"8C", x"8C", x"88", x"44", x"68", x"88", x"88", x"88", x"68", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"89", x"8D", x"8D", x"8D", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"40", x"FF", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"40", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"64", x"64", x"64", x"68", x"88", x"8D", x"8D", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"64", x"68", x"68", x"88", x"88", x"8C", x"8C", x"88", x"44", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"88", x"88", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"88", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"44", x"44", x"24", x"68", x"69", x"44", x"FF", x"00", x"00"),
(x"00", x"00", x"00", x"FF", x"40", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"64", x"64", x"64", x"68", x"88", x"8C", x"AD", x"88", x"68", x"68", x"68", x"64", x"64", x"64", x"44", x"44", x"44", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8D", x"8D", x"8D", x"89", x"8D", x"8C", x"88", x"88", x"88", x"68", x"68", x"68", x"88", x"88", x"88", x"8C", x"8C", x"88", x"88", x"68", x"68", x"44", x"44", x"44", x"00", x"6E", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"B2", x"00", x"68", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"68", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"88", x"89", x"8C", x"88", x"68", x"64", x"44", x"20", x"20", x"44", x"44", x"44", x"68", x"8D", x"6D", x"FF", x"00", x"00", x"00"),
(x"00", x"00", x"FF", x"68", x"89", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"44", x"40", x"44", x"88", x"88", x"68", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"44", x"64", x"68", x"88", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"8D", x"8D", x"8D", x"8C", x"88", x"88", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"88", x"88", x"68", x"88", x"88", x"88", x"88", x"68", x"68", x"6D", x"69", x"FF", x"00", x"00", x"00"),
(x"00", x"00", x"FF", x"64", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"44", x"64", x"64", x"64", x"44", x"44", x"44", x"40", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"44", x"44", x"68", x"88", x"88", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8C", x"88", x"8C", x"88", x"88", x"88", x"88", x"88", x"68", x"64", x"68", x"68", x"69", x"68", x"FF", x"00", x"00", x"00"),
(x"00", x"00", x"B2", x"DB", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"64", x"64", x"64", x"68", x"64", x"64", x"64", x"68", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"44", x"44", x"40", x"20", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"64", x"64", x"64", x"68", x"64", x"44", x"44", x"44", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"64", x"44", x"44", x"44", x"68", x"48", x"FF", x"00", x"00", x"00"),
(x"00", x"00", x"6D", x"40", x"64", x"64", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"64", x"68", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"44", x"44", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"44", x"44", x"44", x"44", x"44", x"64", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"20", x"44", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"64", x"44", x"44", x"44", x"44", x"68", x"44", x"FF", x"00", x"00", x"00"),
(x"00", x"FF", x"88", x"8D", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"44", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"44", x"44", x"44", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"64", x"44", x"44", x"44", x"44", x"69", x"44", x"FF", x"00", x"00", x"00"),
(x"00", x"FF", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"68", x"64", x"68", x"68", x"64", x"68", x"68", x"64", x"64", x"64", x"44", x"44", x"64", x"64", x"64", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"64", x"44", x"44", x"44", x"FF", x"00", x"00", x"00"),
(x"00", x"FF", x"64", x"68", x"68", x"44", x"64", x"64", x"64", x"64", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"44", x"44", x"44", x"64", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"44", x"48", x"44", x"FF", x"00", x"00", x"00"),
(x"00", x"FF", x"44", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"44", x"68", x"64", x"44", x"64", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"64", x"64", x"44", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"64", x"64", x"64", x"44", x"44", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"88", x"88", x"68", x"68", x"48", x"44", x"FF", x"00", x"00", x"00"),
(x"00", x"FF", x"44", x"68", x"68", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"8D", x"8D", x"B2", x"DA", x"B1", x"89", x"68", x"68", x"68", x"68", x"68", x"68", x"64", x"64", x"64", x"68", x"64", x"44", x"64", x"64", x"64", x"68", x"68", x"64", x"44", x"44", x"44", x"64", x"64", x"44", x"68", x"89", x"68", x"68", x"68", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"44", x"64", x"64", x"44", x"44", x"44", x"44", x"64", x"68", x"68", x"68", x"68", x"88", x"89", x"8D", x"91", x"92", x"92", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"FF", x"64", x"68", x"68", x"68", x"68", x"64", x"68", x"68", x"68", x"89", x"89", x"68", x"68", x"68", x"89", x"88", x"8D", x"D2", x"FF", x"FF", x"44", x"FF", x"B1", x"88", x"88", x"88", x"89", x"68", x"64", x"68", x"89", x"8D", x"8D", x"89", x"AD", x"B1", x"DA", x"D6", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DA", x"DB", x"8D", x"69", x"89", x"8D", x"8D", x"68", x"69", x"48", x"69", x"69", x"69", x"69", x"68", x"69", x"69", x"69", x"91", x"B6", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000001111110000000000000001111111111111100000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000001111111111111111011111111111111111111111111000000000000011110000000111111100000"),
("0000000011000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("0001111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111110000000"),
("0001111111111111111100011111111111111110000000000000000000000000000001100000000000011111111111111111100000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;
  end process;
end behav;		

--generated with PNGtoVHDL tool by Ben Wellingstein
