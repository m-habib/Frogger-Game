--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity LoseTable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(12 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end LoseTable;

architecture arch of LoseTable is
constant array_size 			: integer := 4288 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal Lose_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  LoseTable_proc: process(resetN, CLK)
    constant Lose_table : table_type := (
---start 0 v

X"E5A2",
X"E813",
X"EB7E",
X"EC78",
X"F060",
X"F060",
X"F34E",
X"F4C5",
X"F6B9",
X"F8AD",
X"FA24",
X"FC18",
X"FD8F",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"04E2",
X"05DC",
X"0753",
X"084D",
X"0947",
X"0A41",
X"0B3B",
X"0C35",
X"0D2F",
X"0EA6",
X"109A",
X"128E",
X"1482",
X"1676",
X"186A",
X"1A5E",
X"1C52",
X"1DC9",
X"1FBD",
X"2134",
X"222E",
X"23A5",
X"249F",
X"251C",
X"2616",
X"2693",
X"2710",
X"278D",
X"280A",
X"280A",
X"2887",
X"2904",
X"2981",
X"2A7B",
X"2AF8",
X"2B75",
X"2BF2",
X"2C6F",
X"2D69",
X"2DE6",
X"2E63",
X"2EE0",
X"2EE0",
X"2F5D",
X"2FDA",
X"3057",
X"3057",
X"30D4",
X"30D4",
X"3151",
X"31CE",
X"324B",
X"324B",
X"324B",
X"324B",
X"324B",
X"324B",
X"324B",
X"32C8",
X"33C2",
X"34BC",
X"3539",
X"35B6",
X"35B6",
X"35B6",
X"35B6",
X"3633",
X"36B0",
X"36B0",
X"3633",
X"3633",
X"3633",
X"372D",
X"3827",
X"38A4",
X"38A4",
X"3827",
X"3827",
X"37AA",
X"37AA",
X"372D",
X"372D",
X"372D",
X"36B0",
X"36B0",
X"3633",
X"3633",
X"35B6",
X"35B6",
X"35B6",
X"35B6",
X"35B6",
X"3539",
X"3539",
X"34BC",
X"343F",
X"33C2",
X"32C8",
X"3151",
X"2FDA",
X"2DE6",
X"2B75",
X"2981",
X"278D",
X"2693",
X"2693",
X"278D",
X"2887",
X"29FE",
X"2AF8",
X"2B75",
X"2AF8",
X"2AF8",
X"2A7B",
X"2A7B",
X"2A7B",
X"2981",
X"280A",
X"251C",
X"222E",
X"1E46",
X"1ADB",
X"1770",
X"1482",
X"1211",
X"101D",
X"0E29",
X"0D2F",
X"0CB2",
X"0CB2",
X"0C35",
X"0C35",
X"0B3B",
X"0A41",
X"084D",
X"055F",
X"02EE",
X"007D",
X"FE89",
X"FC95",
X"FAA1",
X"F92A",
X"F830",
X"F6B9",
X"F542",
X"F448",
X"F2D1",
X"F15A",
X"EFE3",
X"EDEF",
X"EC78",
X"EB7E",
X"EA84",
X"EA07",
X"E90D",
X"E890",
X"E813",
X"E796",
X"E796",
X"E719",
X"E69C",
X"E5A2",
X"E4A8",
X"E3AE",
X"E2B4",
X"E237",
X"E1BA",
X"E13D",
X"E043",
X"DF49",
X"DE4F",
X"DD55",
X"DC5B",
X"DBDE",
X"DB61",
X"DAE4",
X"DA67",
X"D9EA",
X"D8F0",
X"D873",
X"D7F6",
X"D779",
X"D6FC",
X"D67F",
X"D602",
X"D585",
X"D508",
X"D508",
X"D48B",
X"D40E",
X"D391",
X"D314",
X"D297",
X"D297",
X"D21A",
X"D19D",
X"D19D",
X"D120",
X"D0A3",
X"D0A3",
X"D026",
X"D026",
X"CFA9",
X"CFA9",
X"CF2C",
X"CF2C",
X"CF2C",
X"CEAF",
X"CEAF",
X"CE32",
X"CE32",
X"CDB5",
X"CDB5",
X"CDB5",
X"CDB5",
X"CD38",
X"CD38",
X"CD38",
X"CCBB",
X"CCBB",
X"CCBB",
X"CCBB",
X"CCBB",
X"CCBB",
X"CCBB",
X"CCBB",
X"CD38",
X"CD38",
X"CD38",
X"CD38",
X"CDB5",
X"CDB5",
X"CDB5",
X"CE32",
X"CEAF",
X"CF2C",
X"CFA9",
X"D026",
X"D026",
X"D026",
X"D026",
X"D026",
X"D026",
X"D0A3",
X"D0A3",
X"D120",
X"D120",
X"D19D",
X"D19D",
X"D21A",
X"D314",
X"D40E",
X"D48B",
X"D508",
X"D508",
X"D585",
X"D67F",
X"D779",
X"D7F6",
X"D8F0",
X"D9EA",
X"DA67",
X"DA67",
X"DAE4",
X"DB61",
X"DBDE",
X"DC5B",
X"DD55",
X"DE4F",
X"DECC",
X"DFC6",
X"E043",
X"E0C0",
X"E0C0",
X"E1BA",
X"E2B4",
X"E3AE",
X"E4A8",
X"E61F",
X"E719",
X"E813",
X"E98A",
X"EA84",
X"EB01",
X"EBFB",
X"EBFB",
X"EC78",
X"ECF5",
X"ED72",
X"EDEF",
X"EEE9",
X"EFE3",
X"F15A",
X"F2D1",
X"F3CB",
X"F542",
X"F63C",
X"F7B3",
X"F8AD",
X"F92A",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"0000",
X"00FA",
X"01F4",
X"036B",
X"0465",
X"055F",
X"0659",
X"06D6",
X"07D0",
X"084D",
X"08CA",
X"08CA",
X"0947",
X"09C4",
X"0ABE",
X"0BB8",
X"0CB2",
X"0E29",
X"0F23",
X"109A",
X"1194",
X"128E",
X"1388",
X"1405",
X"1482",
X"14FF",
X"15F9",
X"1676",
X"1770",
X"17ED",
X"18E7",
X"1964",
X"1A5E",
X"1ADB",
X"1BD5",
X"1CCF",
X"1D4C",
X"1DC9",
X"1EC3",
X"1F40",
X"1FBD",
X"203A",
X"20B7",
X"2134",
X"21B1",
X"222E",
X"22AB",
X"22AB",
X"2328",
X"23A5",
X"23A5",
X"2422",
X"249F",
X"251C",
X"2599",
X"2599",
X"2616",
X"2693",
X"2710",
X"2710",
X"278D",
X"278D",
X"280A",
X"280A",
X"280A",
X"278D",
X"278D",
X"278D",
X"278D",
X"278D",
X"280A",
X"280A",
X"280A",
X"2887",
X"2887",
X"2887",
X"2887",
X"2904",
X"2904",
X"2904",
X"2904",
X"2887",
X"2887",
X"2904",
X"2904",
X"2904",
X"2904",
X"2904",
X"2904",
X"2887",
X"2887",
X"2887",
X"2887",
X"2887",
X"280A",
X"280A",
X"280A",
X"280A",
X"278D",
X"278D",
X"278D",
X"2710",
X"2710",
X"2710",
X"2693",
X"2693",
X"2693",
X"2616",
X"2616",
X"2616",
X"2599",
X"2599",
X"2599",
X"251C",
X"251C",
X"251C",
X"249F",
X"249F",
X"249F",
X"2422",
X"2422",
X"23A5",
X"23A5",
X"2328",
X"2328",
X"2328",
X"22AB",
X"22AB",
X"222E",
X"222E",
X"21B1",
X"21B1",
X"2134",
X"20B7",
X"20B7",
X"203A",
X"203A",
X"1FBD",
X"1FBD",
X"1F40",
X"1EC3",
X"1E46",
X"1DC9",
X"1D4C",
X"1CCF",
X"1C52",
X"1BD5",
X"1B58",
X"1ADB",
X"1A5E",
X"19E1",
X"1964",
X"18E7",
X"186A",
X"17ED",
X"17ED",
X"1770",
X"16F3",
X"16F3",
X"1676",
X"1676",
X"15F9",
X"157C",
X"14FF",
X"1405",
X"1388",
X"128E",
X"128E",
X"1211",
X"1194",
X"1194",
X"1117",
X"109A",
X"109A",
X"101D",
X"0FA0",
X"0F23",
X"0EA6",
X"0E29",
X"0DAC",
X"0D2F",
X"0CB2",
X"0C35",
X"0B3B",
X"0ABE",
X"0A41",
X"09C4",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"0753",
X"06D6",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"04E2",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FF06",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"F9A7",
X"F8AD",
X"F7B3",
X"F6B9",
X"F63C",
X"F542",
X"F4C5",
X"F448",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F34E",
X"F34E",
X"F2D1",
X"F254",
X"F15A",
X"F060",
X"EF66",
X"EEE9",
X"EE6C",
X"EE6C",
X"EE6C",
X"EDEF",
X"EDEF",
X"EDEF",
X"ED72",
X"ED72",
X"ECF5",
X"ECF5",
X"EC78",
X"EBFB",
X"EBFB",
X"EB7E",
X"EB7E",
X"EB01",
X"EA84",
X"EA84",
X"EA07",
X"EA07",
X"E98A",
X"E98A",
X"E90D",
X"E90D",
X"E890",
X"E890",
X"E813",
X"E813",
X"E796",
X"E796",
X"E719",
X"E719",
X"E69C",
X"E69C",
X"E69C",
X"E61F",
X"E61F",
X"E61F",
X"E5A2",
X"E5A2",
X"E525",
X"E525",
X"E4A8",
X"E42B",
X"E42B",
X"E3AE",
X"E3AE",
X"E3AE",
X"E331",
X"E331",
X"E331",
X"E331",
X"E2B4",
X"E2B4",
X"E2B4",
X"E237",
X"E237",
X"E237",
X"E237",
X"E1BA",
X"E1BA",
X"E1BA",
X"E13D",
X"E13D",
X"E13D",
X"E0C0",
X"E0C0",
X"E043",
X"E043",
X"DFC6",
X"DFC6",
X"DFC6",
X"DF49",
X"DF49",
X"DF49",
X"DF49",
X"DECC",
X"DECC",
X"DECC",
X"DE4F",
X"DE4F",
X"DE4F",
X"DDD2",
X"DDD2",
X"DE4F",
X"DE4F",
X"DECC",
X"DECC",
X"DECC",
X"DECC",
X"DE4F",
X"DE4F",
X"DDD2",
X"DDD2",
X"DDD2",
X"DDD2",
X"DDD2",
X"DDD2",
X"DDD2",
X"DDD2",
X"DDD2",
X"DE4F",
X"DECC",
X"DF49",
X"DF49",
X"DFC6",
X"DFC6",
X"E043",
X"E0C0",
X"E0C0",
X"E13D",
X"E1BA",
X"E1BA",
X"E237",
X"E2B4",
X"E331",
X"E331",
X"E3AE",
X"E42B",
X"E4A8",
X"E525",
X"E5A2",
X"E5A2",
X"E61F",
X"E719",
X"E796",
X"E796",
X"E813",
X"E813",
X"E813",
X"E890",
X"E890",
X"E890",
X"E890",
X"E90D",
X"E98A",
X"EA84",
X"EB01",
X"EBFB",
X"EC78",
X"ED72",
X"EDEF",
X"EE6C",
X"EE6C",
X"EE6C",
X"EE6C",
X"EE6C",
X"EE6C",
X"EEE9",
X"EEE9",
X"EF66",
X"EFE3",
X"F060",
X"F0DD",
X"F1D7",
X"F2D1",
X"F34E",
X"F448",
X"F4C5",
X"F5BF",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"05DC",
X"0659",
X"06D6",
X"07D0",
X"084D",
X"08CA",
X"0947",
X"0947",
X"09C4",
X"09C4",
X"0A41",
X"0A41",
X"0A41",
X"0ABE",
X"0B3B",
X"0BB8",
X"0C35",
X"0CB2",
X"0D2F",
X"0DAC",
X"0E29",
X"0EA6",
X"0EA6",
X"0F23",
X"0FA0",
X"0FA0",
X"101D",
X"101D",
X"101D",
X"109A",
X"109A",
X"1117",
X"1117",
X"1194",
X"1194",
X"1211",
X"1211",
X"128E",
X"128E",
X"130B",
X"130B",
X"1388",
X"1388",
X"1405",
X"1405",
X"1405",
X"1482",
X"1482",
X"1482",
X"1482",
X"1482",
X"1482",
X"14FF",
X"14FF",
X"14FF",
X"14FF",
X"14FF",
X"14FF",
X"14FF",
X"14FF",
X"157C",
X"157C",
X"157C",
X"157C",
X"15F9",
X"15F9",
X"15F9",
X"15F9",
X"1676",
X"1676",
X"1676",
X"1676",
X"1676",
X"1676",
X"1676",
X"16F3",
X"16F3",
X"16F3",
X"16F3",
X"16F3",
X"16F3",
X"1770",
X"1770",
X"1770",
X"1770",
X"1770",
X"17ED",
X"17ED",
X"17ED",
X"17ED",
X"17ED",
X"17ED",
X"186A",
X"186A",
X"186A",
X"186A",
X"186A",
X"186A",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"1964",
X"1964",
X"1964",
X"1964",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"1964",
X"1964",
X"1964",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"19E1",
X"1964",
X"1964",
X"1964",
X"1964",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"18E7",
X"186A",
X"186A",
X"17ED",
X"17ED",
X"1770",
X"16F3",
X"16F3",
X"1676",
X"1676",
X"15F9",
X"15F9",
X"157C",
X"14FF",
X"14FF",
X"1482",
X"1405",
X"1388",
X"1388",
X"130B",
X"130B",
X"128E",
X"128E",
X"128E",
X"128E",
X"1211",
X"1211",
X"1211",
X"1194",
X"1117",
X"1117",
X"109A",
X"101D",
X"0FA0",
X"0EA6",
X"0E29",
X"0DAC",
X"0DAC",
X"0D2F",
X"0D2F",
X"0CB2",
X"0CB2",
X"0C35",
X"0C35",
X"0BB8",
X"0B3B",
X"0ABE",
X"0A41",
X"09C4",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"0753",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F5BF",
X"F542",
X"F4C5",
X"F4C5",
X"F448",
X"F3CB",
X"F3CB",
X"F34E",
X"F2D1",
X"F2D1",
X"F2D1",
X"F254",
X"F254",
X"F1D7",
X"F1D7",
X"F15A",
X"F15A",
X"F0DD",
X"F060",
X"F060",
X"EFE3",
X"EFE3",
X"EF66",
X"EF66",
X"EF66",
X"EF66",
X"EF66",
X"EF66",
X"EF66",
X"EF66",
X"EF66",
X"EF66",
X"EEE9",
X"EEE9",
X"EEE9",
X"EE6C",
X"EE6C",
X"EDEF",
X"EDEF",
X"EDEF",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"EC78",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ECF5",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"ED72",
X"EDEF",
X"EDEF",
X"EDEF",
X"EE6C",
X"EE6C",
X"EE6C",
X"EEE9",
X"EEE9",
X"EF66",
X"EFE3",
X"EFE3",
X"F060",
X"F060",
X"F0DD",
X"F0DD",
X"F0DD",
X"F0DD",
X"F0DD",
X"F15A",
X"F15A",
X"F1D7",
X"F1D7",
X"F254",
X"F254",
X"F2D1",
X"F34E",
X"F34E",
X"F3CB",
X"F3CB",
X"F448",
X"F448",
X"F4C5",
X"F4C5",
X"F542",
X"F5BF",
X"F5BF",
X"F63C",
X"F63C",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F7B3",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"FAA1",
X"FB1E",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"0947",
X"09C4",
X"09C4",
X"0A41",
X"0A41",
X"0ABE",
X"0ABE",
X"0ABE",
X"0ABE",
X"0ABE",
X"0B3B",
X"0B3B",
X"0B3B",
X"0B3B",
X"0B3B",
X"0B3B",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0C35",
X"0C35",
X"0C35",
X"0CB2",
X"0CB2",
X"0CB2",
X"0D2F",
X"0D2F",
X"0D2F",
X"0DAC",
X"0DAC",
X"0E29",
X"0E29",
X"0E29",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0EA6",
X"0F23",
X"0F23",
X"0F23",
X"0FA0",
X"0FA0",
X"0FA0",
X"101D",
X"101D",
X"101D",
X"101D",
X"101D",
X"109A",
X"109A",
X"109A",
X"109A",
X"109A",
X"109A",
X"109A",
X"109A",
X"109A",
X"109A",
X"109A",
X"1117",
X"1117",
X"1117",
X"1194",
X"1194",
X"1211",
X"128E",
X"128E",
X"128E",
X"128E",
X"128E",
X"128E",
X"1211",
X"1211",
X"1211",
X"1211",
X"1194",
X"1194",
X"1194",
X"1194",
X"1194",
X"1194",
X"1211",
X"1211",
X"1211",
X"1211",
X"1194",
X"1194",
X"1194",
X"1194",
X"1194",
X"1194",
X"1117",
X"1117",
X"1117",
X"109A",
X"109A",
X"109A",
X"101D",
X"101D",
X"0FA0",
X"0FA0",
X"0F23",
X"0F23",
X"0EA6",
X"0EA6",
X"0EA6",
X"0E29",
X"0E29",
X"0E29",
X"0E29",
X"0DAC",
X"0DAC",
X"0D2F",
X"0D2F",
X"0CB2",
X"0C35",
X"0BB8",
X"0BB8",
X"0B3B",
X"0ABE",
X"0A41",
X"09C4",
X"0947",
X"08CA",
X"08CA",
X"084D",
X"07D0",
X"0753",
X"0753",
X"06D6",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F736",
X"F736",
X"F736",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F5BF",
X"F5BF",
X"F5BF",
X"F5BF",
X"F5BF",
X"F542",
X"F542",
X"F542",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F4C5",
X"F4C5",
X"F542",
X"F542",
X"F542",
X"F5BF",
X"F5BF",
X"F5BF",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"07D0",
X"07D0",
X"07D0",
X"07D0",
X"0753",
X"0753",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"0659",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F63C",
X"F63C",
X"F63C",
X"F5BF",
X"F5BF",
X"F5BF",
X"F542",
X"F542",
X"F542",
X"F542",
X"F4C5",
X"F4C5",
X"F448",
X"F448",
X"F448",
X"F448",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F34E",
X"F34E",
X"F34E",
X"F2D1",
X"F2D1",
X"F2D1",
X"F2D1",
X"F254",
X"F254",
X"F254",
X"F1D7",
X"F1D7",
X"F1D7",
X"F1D7",
X"F1D7",
X"F1D7",
X"F1D7",
X"F1D7",
X"F1D7",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F1D7",
X"F1D7",
X"F1D7",
X"F1D7",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F15A",
X"F1D7",
X"F1D7",
X"F1D7",
X"F254",
X"F254",
X"F254",
X"F2D1",
X"F2D1",
X"F2D1",
X"F34E",
X"F34E",
X"F3CB",
X"F3CB",
X"F3CB",
X"F3CB",
X"F448",
X"F448",
X"F448",
X"F448",
X"F4C5",
X"F4C5",
X"F542",
X"F542",
X"F542",
X"F5BF",
X"F5BF",
X"F5BF",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F736",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"0947",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0ABE",
X"0ABE",
X"0ABE",
X"0B3B",
X"0B3B",
X"0B3B",
X"0B3B",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0C35",
X"0C35",
X"0C35",
X"0C35",
X"0C35",
X"0C35",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0D2F",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0CB2",
X"0C35",
X"0C35",
X"0C35",
X"0C35",
X"0C35",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0BB8",
X"0B3B",
X"0B3B",
X"0ABE",
X"0ABE",
X"0ABE",
X"0A41",
X"0A41",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"0947",
X"0947",
X"0947",
X"0947",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"084D",
X"084D",
X"084D",
X"07D0",
X"07D0",
X"0753",
X"0753",
X"06D6",
X"06D6",
X"0659",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"0947",
X"0947",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0ABE",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"0A41",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"09C4",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"0947",
X"08CA",
X"08CA",
X"08CA",
X"08CA",
X"084D",
X"084D",
X"084D",
X"07D0",
X"07D0",
X"07D0",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"F92A",
X"F92A",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F830",
X"F830",
X"F830",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F736",
X"F736",
X"F736",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F63C",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F6B9",
X"F736",
X"F736",
X"F736",
X"F736",
X"F7B3",
X"F7B3",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F830",
X"F830",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"055F",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"07D0",
X"07D0",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"084D",
X"07D0",
X"07D0",
X"07D0",
X"07D0",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"0753",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"0659",
X"0659",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000"




 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= Lose_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;