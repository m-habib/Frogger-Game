--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity JumpTable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(11 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end JumpTable;

architecture arch of JumpTable is
constant array_size 			: integer := 3528 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal Jump_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  JumpTable_proc: process(resetN, CLK)
    constant Jump_table : table_type := (
---start 0 v

X"0000",
X"01F4",
X"0465",
X"0659",
X"08CA",
X"0ABE",
X"0CB2",
X"0EA6",
X"109A",
X"128E",
X"1405",
X"15F9",
X"1770",
X"18E7",
X"1A5E",
X"1B58",
X"1C52",
X"1D4C",
X"1DC9",
X"1E46",
X"1EC3",
X"1F40",
X"1F40",
X"1F40",
X"1EC3",
X"1E46",
X"1DC9",
X"1D4C",
X"1C52",
X"1B58",
X"1A5E",
X"18E7",
X"1770",
X"15F9",
X"1405",
X"128E",
X"109A",
X"0EA6",
X"0CB2",
X"0A41",
X"084D",
X"0659",
X"03E8",
X"0177",
X"FF83",
X"FD12",
X"FAA1",
X"F8AD",
X"F63C",
X"F448",
X"F1D7",
X"EFE3",
X"EDEF",
X"EBFB",
X"EA84",
X"E890",
X"E719",
X"E5A2",
X"E4A8",
X"E3AE",
X"E2B4",
X"E1BA",
X"E0C0",
X"E043",
X"E043",
X"DFC6",
X"DFC6",
X"E043",
X"E043",
X"E0C0",
X"E1BA",
X"E237",
X"E331",
X"E4A8",
X"E5A2",
X"E719",
X"E890",
X"EA84",
X"EBFB",
X"EDEF",
X"EFE3",
X"F254",
X"F448",
X"F6B9",
X"F8AD",
X"FB1E",
X"FD8F",
X"FF83",
X"01F4",
X"0465",
X"06D6",
X"08CA",
X"0B3B",
X"0D2F",
X"0FA0",
X"1194",
X"1388",
X"14FF",
X"16F3",
X"186A",
X"19E1",
X"1B58",
X"1C52",
X"1D4C",
X"1E46",
X"1EC3",
X"1F40",
X"1FBD",
X"1FBD",
X"1FBD",
X"1FBD",
X"1F40",
X"1EC3",
X"1E46",
X"1D4C",
X"1C52",
X"1B58",
X"19E1",
X"186A",
X"1676",
X"14FF",
X"130B",
X"1117",
X"0F23",
X"0D2F",
X"0ABE",
X"084D",
X"0659",
X"03E8",
X"0177",
X"FF06",
X"FC95",
X"FA24",
X"F7B3",
X"F5BF",
X"F34E",
X"F0DD",
X"EEE9",
X"ECF5",
X"EB01",
X"E90D",
X"E796",
X"E61F",
X"E4A8",
X"E331",
X"E237",
X"E13D",
X"E043",
X"DFC6",
X"DF49",
X"DF49",
X"DF49",
X"DF49",
X"DFC6",
X"E043",
X"E0C0",
X"E1BA",
X"E2B4",
X"E3AE",
X"E525",
X"E69C",
X"E813",
X"EA07",
X"EBFB",
X"EDEF",
X"EFE3",
X"F1D7",
X"F448",
X"F6B9",
X"F92A",
X"FB9B",
X"FE0C",
X"007D",
X"02EE",
X"055F",
X"07D0",
X"0A41",
X"0C35",
X"0EA6",
X"109A",
X"130B",
X"14FF",
X"1676",
X"186A",
X"19E1",
X"1B58",
X"1CCF",
X"1DC9",
X"1EC3",
X"1F40",
X"203A",
X"203A",
X"20B7",
X"20B7",
X"20B7",
X"203A",
X"1FBD",
X"1EC3",
X"1E46",
X"1CCF",
X"1BD5",
X"1A5E",
X"18E7",
X"16F3",
X"14FF",
X"130B",
X"1117",
X"0F23",
X"0CB2",
X"0A41",
X"07D0",
X"055F",
X"02EE",
X"007D",
X"FE0C",
X"FB9B",
X"F92A",
X"F6B9",
X"F448",
X"F1D7",
X"EF66",
X"ED72",
X"EB7E",
X"E98A",
X"E796",
X"E5A2",
X"E42B",
X"E331",
X"E1BA",
X"E0C0",
X"DFC6",
X"DF49",
X"DECC",
X"DE4F",
X"DE4F",
X"DECC",
X"DECC",
X"DF49",
X"E043",
X"E0C0",
X"E237",
X"E331",
X"E4A8",
X"E61F",
X"E813",
X"EA07",
X"EBFB",
X"EDEF",
X"F060",
X"F254",
X"F4C5",
X"F736",
X"F9A7",
X"FC95",
X"FF06",
X"0177",
X"03E8",
X"06D6",
X"0947",
X"0BB8",
X"0E29",
X"101D",
X"128E",
X"1482",
X"1676",
X"186A",
X"1A5E",
X"1BD5",
X"1D4C",
X"1E46",
X"1F40",
X"203A",
X"20B7",
X"2134",
X"2134",
X"2134",
X"2134",
X"20B7",
X"203A",
X"1FBD",
X"1EC3",
X"1D4C",
X"1C52",
X"1A5E",
X"18E7",
X"16F3",
X"14FF",
X"130B",
X"109A",
X"0EA6",
X"0C35",
X"09C4",
X"06D6",
X"0465",
X"01F4",
X"FF06",
X"FC95",
X"FA24",
X"F736",
X"F4C5",
X"F254",
X"EFE3",
X"ED72",
X"EB7E",
X"E98A",
X"E796",
X"E5A2",
X"E42B",
X"E2B4",
X"E13D",
X"E043",
X"DF49",
X"DECC",
X"DE4F",
X"DDD2",
X"DDD2",
X"DDD2",
X"DE4F",
X"DECC",
X"DF49",
X"E043",
X"E1BA",
X"E2B4",
X"E4A8",
X"E61F",
X"E813",
X"EA07",
X"EBFB",
X"EE6C",
X"F0DD",
X"F34E",
X"F5BF",
X"F830",
X"FB1E",
X"FD8F",
X"007D",
X"02EE",
X"05DC",
X"084D",
X"0ABE",
X"0DAC",
X"101D",
X"1211",
X"1482",
X"1676",
X"186A",
X"1A5E",
X"1BD5",
X"1D4C",
X"1EC3",
X"1FBD",
X"20B7",
X"2134",
X"21B1",
X"222E",
X"222E",
X"222E",
X"21B1",
X"20B7",
X"203A",
X"1F40",
X"1DC9",
X"1C52",
X"1ADB",
X"18E7",
X"16F3",
X"14FF",
X"128E",
X"109A",
X"0DAC",
X"0B3B",
X"08CA",
X"05DC",
X"036B",
X"007D",
X"FD8F",
X"FB1E",
X"F830",
X"F5BF",
X"F2D1",
X"F060",
X"EDEF",
X"EB7E",
X"E98A",
X"E796",
X"E5A2",
X"E3AE",
X"E237",
X"E0C0",
X"DFC6",
X"DECC",
X"DDD2",
X"DD55",
X"DD55",
X"DCD8",
X"DD55",
X"DD55",
X"DE4F",
X"DECC",
X"DFC6",
X"E13D",
X"E2B4",
X"E42B",
X"E61F",
X"E813",
X"EA07",
X"EC78",
X"EEE9",
X"F15A",
X"F3CB",
X"F6B9",
X"F92A",
X"FC18",
X"FF06",
X"01F4",
X"0465",
X"0753",
X"0A41",
X"0CB2",
X"0F23",
X"1211",
X"1405",
X"1676",
X"186A",
X"1A5E",
X"1C52",
X"1DC9",
X"1F40",
X"203A",
X"2134",
X"222E",
X"22AB",
X"22AB",
X"22AB",
X"22AB",
X"222E",
X"21B1",
X"20B7",
X"1FBD",
X"1E46",
X"1CCF",
X"1ADB",
X"18E7",
X"16F3",
X"14FF",
X"128E",
X"101D",
X"0D2F",
X"0ABE",
X"07D0",
X"04E2",
X"01F4",
X"FF83",
X"FC95",
X"F9A7",
X"F6B9",
X"F3CB",
X"F15A",
X"EEE9",
X"EBFB",
X"EA07",
X"E796",
X"E5A2",
X"E3AE",
X"E237",
X"E0C0",
X"DF49",
X"DE4F",
X"DD55",
X"DCD8",
X"DC5B",
X"DC5B",
X"DC5B",
X"DCD8",
X"DD55",
X"DE4F",
X"DF49",
X"E0C0",
X"E237",
X"E3AE",
X"E5A2",
X"E796",
X"EA07",
X"EC78",
X"EEE9",
X"F1D7",
X"F448",
X"F736",
X"FA24",
X"FD12",
X"0000",
X"02EE",
X"05DC",
X"08CA",
X"0BB8",
X"0E29",
X"1117",
X"1388",
X"15F9",
X"17ED",
X"1A5E",
X"1C52",
X"1DC9",
X"1F40",
X"20B7",
X"21B1",
X"22AB",
X"2328",
X"23A5",
X"23A5",
X"2328",
X"2328",
X"222E",
X"2134",
X"203A",
X"1EC3",
X"1D4C",
X"1B58",
X"1964",
X"1770",
X"14FF",
X"128E",
X"101D",
X"0D2F",
X"0A41",
X"0753",
X"0465",
X"0177",
X"FE89",
X"FB9B",
X"F8AD",
X"F5BF",
X"F2D1",
X"EFE3",
X"ED72",
X"EA84",
X"E890",
X"E61F",
X"E42B",
X"E237",
X"E0C0",
X"DF49",
X"DDD2",
X"DCD8",
X"DC5B",
X"DBDE",
X"DBDE",
X"DBDE",
X"DBDE",
X"DCD8",
X"DD55",
X"DE4F",
X"DFC6",
X"E13D",
X"E331",
X"E525",
X"E719",
X"E98A",
X"EBFB",
X"EEE9",
X"F15A",
X"F448",
X"F736",
X"FA24",
X"FD8F",
X"007D",
X"036B",
X"0659",
X"09C4",
X"0CB2",
X"0F23",
X"1211",
X"1482",
X"16F3",
X"1964",
X"1B58",
X"1D4C",
X"1F40",
X"20B7",
X"21B1",
X"22AB",
X"23A5",
X"2422",
X"2422",
X"2422",
X"23A5",
X"2328",
X"222E",
X"2134",
X"1FBD",
X"1E46",
X"1C52",
X"1A5E",
X"186A",
X"15F9",
X"130B",
X"109A",
X"0DAC",
X"0ABE",
X"07D0",
X"04E2",
X"0177",
X"FE89",
X"FB1E",
X"F830",
X"F542",
X"F254",
X"EF66",
X"EC78",
X"EA07",
X"E796",
X"E525",
X"E331",
X"E13D",
X"DFC6",
X"DE4F",
X"DCD8",
X"DC5B",
X"DB61",
X"DAE4",
X"DAE4",
X"DB61",
X"DBDE",
X"DC5B",
X"DD55",
X"DECC",
X"E043",
X"E1BA",
X"E3AE",
X"E61F",
X"E890",
X"EB01",
X"ED72",
X"F060",
X"F34E",
X"F63C",
X"F9A7",
X"FC95",
X"0000",
X"02EE",
X"0659",
X"0947",
X"0CB2",
X"0FA0",
X"128E",
X"14FF",
X"1770",
X"19E1",
X"1C52",
X"1E46",
X"1FBD",
X"2134",
X"22AB",
X"23A5",
X"2422",
X"249F",
X"249F",
X"249F",
X"2422",
X"23A5",
X"22AB",
X"2134",
X"1FBD",
X"1E46",
X"1C52",
X"19E1",
X"1770",
X"14FF",
X"1211",
X"0F23",
X"0C35",
X"0947",
X"05DC",
X"0271",
X"FF83",
X"FC18",
X"F8AD",
X"F5BF",
X"F2D1",
X"EF66",
X"EC78",
X"EA07",
X"E796",
X"E525",
X"E2B4",
X"E0C0",
X"DF49",
X"DDD2",
X"DC5B",
X"DB61",
X"DAE4",
X"DA67",
X"DA67",
X"DA67",
X"DAE4",
X"DBDE",
X"DCD8",
X"DE4F",
X"DFC6",
X"E1BA",
X"E3AE",
X"E61F",
X"E890",
X"EB7E",
X"EE6C",
X"F15A",
X"F448",
X"F7B3",
X"FB1E",
X"FE0C",
X"0177",
X"04E2",
X"084D",
X"0B3B",
X"0EA6",
X"1194",
X"1482",
X"16F3",
X"19E1",
X"1BD5",
X"1E46",
X"1FBD",
X"21B1",
X"2328",
X"2422",
X"249F",
X"251C",
X"2599",
X"251C",
X"251C",
X"2422",
X"2328",
X"21B1",
X"203A",
X"1EC3",
X"1C52",
X"1A5E",
X"1770",
X"14FF",
X"1211",
X"0F23",
X"0BB8",
X"08CA",
X"055F",
X"01F4",
X"FE89",
X"FB1E",
X"F7B3",
X"F448",
X"F15A",
X"EDEF",
X"EB01",
X"E890",
X"E5A2",
X"E331",
X"E13D",
X"DF49",
X"DDD2",
X"DC5B",
X"DB61",
X"DA67",
X"D9EA",
X"D9EA",
X"D9EA",
X"DA67",
X"DAE4",
X"DBDE",
X"DD55",
X"DF49",
X"E0C0",
X"E331",
X"E5A2",
X"E813",
X"EB01",
X"EDEF",
X"F0DD",
X"F448",
X"F7B3",
X"FB1E",
X"FE89",
X"01F4",
X"055F",
X"08CA",
X"0C35",
X"0F23",
X"128E",
X"157C",
X"17ED",
X"1ADB",
X"1CCF",
X"1F40",
X"2134",
X"22AB",
X"2422",
X"251C",
X"2599",
X"2616",
X"2616",
X"2599",
X"251C",
X"2422",
X"2328",
X"21B1",
X"1FBD",
X"1DC9",
X"1B58",
X"18E7",
X"1676",
X"1388",
X"101D",
X"0D2F",
X"09C4",
X"0659",
X"0271",
X"FF06",
X"FB9B",
X"F830",
X"F4C5",
X"F15A",
X"EDEF",
X"EB01",
X"E813",
X"E5A2",
X"E331",
X"E0C0",
X"DECC",
X"DCD8",
X"DBDE",
X"DA67",
X"D9EA",
X"D96D",
X"D8F0",
X"D96D",
X"D9EA",
X"DAE4",
X"DBDE",
X"DD55",
X"DF49",
X"E13D",
X"E331",
X"E61F",
X"E890",
X"EB7E",
X"EEE9",
X"F254",
X"F5BF",
X"F92A",
X"FC95",
X"0000",
X"03E8",
X"0753",
X"0ABE",
X"0E29",
X"1194",
X"1482",
X"1770",
X"1A5E",
X"1CCF",
X"1F40",
X"2134",
X"22AB",
X"2422",
X"251C",
X"2616",
X"2693",
X"2693",
X"2693",
X"2616",
X"251C",
X"23A5",
X"222E",
X"203A",
X"1E46",
X"1BD5",
X"1964",
X"1676",
X"130B",
X"101D",
X"0CB2",
X"0947",
X"055F",
X"01F4",
X"FE0C",
X"FAA1",
X"F6B9",
X"F34E",
X"EFE3",
X"EC78",
X"E98A",
X"E69C",
X"E42B",
X"E13D",
X"DF49",
X"DD55",
X"DBDE",
X"DA67",
X"D96D",
X"D8F0",
X"D873",
X"D873",
X"D8F0",
X"D9EA",
X"DAE4",
X"DC5B",
X"DDD2",
X"E043",
X"E237",
X"E525",
X"E813",
X"EB01",
X"EDEF",
X"F15A",
X"F542",
X"F8AD",
X"FC18",
X"0000",
X"03E8",
X"0753",
X"0B3B",
X"0EA6",
X"1211",
X"14FF",
X"186A",
X"1ADB",
X"1DC9",
X"1FBD",
X"222E",
X"23A5",
X"251C",
X"2616",
X"2710",
X"2710",
X"2710",
X"2710",
X"2616",
X"251C",
X"23A5",
X"21B1",
X"1FBD",
X"1DC9",
X"1ADB",
X"17ED",
X"14FF",
X"1194",
X"0E29",
X"0ABE",
X"06D6",
X"036B",
X"FF83",
X"FB9B",
X"F7B3",
X"F448",
X"F0DD",
X"ED72",
X"EA07",
X"E69C",
X"E42B",
X"E13D",
X"DF49",
X"DCD8",
X"DB61",
X"D9EA",
X"D8F0",
X"D873",
X"D7F6",
X"D7F6",
X"D873",
X"D96D",
X"DA67",
X"DBDE",
X"DDD2",
X"DFC6",
X"E237",
X"E525",
X"E813",
X"EB7E",
X"EE6C",
X"F254",
X"F5BF",
X"F9A7",
X"FD8F",
X"0177",
X"055F",
X"08CA",
X"0CB2",
X"101D",
X"1388",
X"16F3",
X"19E1",
X"1CCF",
X"1F40",
X"21B1",
X"23A5",
X"251C",
X"2693",
X"2710",
X"278D",
X"280A",
X"278D",
X"2710",
X"2616",
X"249F",
X"22AB",
X"20B7",
X"1E46",
X"1BD5",
X"18E7",
X"157C",
X"128E",
X"0EA6",
X"0B3B",
X"0753",
X"036B",
X"FF83",
X"FB9B",
X"F7B3",
X"F3CB",
X"F060",
X"EC78",
X"E90D",
X"E61F",
X"E331",
X"E0C0",
X"DE4F",
X"DC5B",
X"DA67",
X"D8F0",
X"D7F6",
X"D779",
X"D779",
X"D779",
X"D7F6",
X"D8F0",
X"DA67",
X"DC5B",
X"DE4F",
X"E0C0",
X"E331",
X"E61F",
X"E98A",
X"ECF5",
X"F060",
X"F448",
X"F830",
X"FC18",
X"0000",
X"03E8",
X"07D0",
X"0BB8",
X"0FA0",
X"130B",
X"1676",
X"19E1",
X"1CCF",
X"1F40",
X"21B1",
X"23A5",
X"2599",
X"2693",
X"278D",
X"280A",
X"2887",
X"280A",
X"278D",
X"2693",
X"251C",
X"2328",
X"2134",
X"1EC3",
X"1BD5",
X"18E7",
X"157C",
X"1211",
X"0E29",
X"0A41",
X"0659",
X"0271",
X"FE89",
X"FA24",
X"F63C",
X"F254",
X"EE6C",
X"EB01",
X"E796",
X"E42B",
X"E1BA",
X"DECC",
X"DCD8",
X"DAE4",
X"D8F0",
X"D7F6",
X"D779",
X"D6FC",
X"D6FC",
X"D779",
X"D873",
X"D96D",
X"DAE4",
X"DD55",
X"DF49",
X"E237",
X"E525",
X"E890",
X"EBFB",
X"EF66",
X"F34E",
X"F736",
X"FB9B",
X"FF83",
X"03E8",
X"07D0",
X"0BB8",
X"0FA0",
X"1388",
X"16F3",
X"1A5E",
X"1D4C",
X"203A",
X"22AB",
X"249F",
X"2616",
X"278D",
X"2887",
X"2904",
X"2904",
X"2887",
X"278D",
X"2693",
X"251C",
X"2328",
X"20B7",
X"1DC9",
X"1ADB",
X"17ED",
X"1405",
X"109A",
X"0CB2",
X"08CA",
X"0465",
X"0000",
X"FC18",
X"F7B3",
X"F3CB",
X"EFE3",
X"EBFB",
X"E890",
X"E525",
X"E237",
X"DF49",
X"DCD8",
X"DAE4",
X"D8F0",
X"D779",
X"D6FC",
X"D67F",
X"D67F",
X"D67F",
X"D779",
X"D8F0",
X"DA67",
X"DC5B",
X"DECC",
X"E1BA",
X"E4A8",
X"E813",
X"EBFB",
X"EF66",
X"F3CB",
X"F7B3",
X"FC18",
X"0000",
X"0465",
X"08CA",
X"0CB2",
X"109A",
X"1482",
X"17ED",
X"1B58",
X"1EC3",
X"2134",
X"23A5",
X"2599",
X"2710",
X"2887",
X"2904",
X"2981",
X"2981",
X"2904",
X"278D",
X"2693",
X"249F",
X"222E",
X"1FBD",
X"1CCF",
X"1964",
X"15F9",
X"1211",
X"0E29",
X"0A41",
X"05DC",
X"0177",
X"FD12",
X"F8AD",
X"F4C5",
X"F060",
X"EC78",
X"E890",
X"E525",
X"E237",
X"DF49",
X"DC5B",
X"DA67",
X"D873",
X"D6FC",
X"D67F",
X"D602",
X"D602",
X"D602",
X"D6FC",
X"D873",
X"DA67",
X"DC5B",
X"DECC",
X"E1BA",
X"E525",
X"E890",
X"EC78",
X"F060",
X"F448",
X"F8AD",
X"FD12",
X"0177",
X"05DC",
X"0A41",
X"0EA6",
X"128E",
X"1676",
X"19E1",
X"1D4C",
X"203A",
X"22AB",
X"251C",
X"2710",
X"2887",
X"2981",
X"29FE",
X"29FE",
X"2981",
X"2887",
X"278D",
X"2599",
X"23A5",
X"20B7",
X"1DC9",
X"1ADB",
X"16F3",
X"130B",
X"0F23",
X"0ABE",
X"0659",
X"01F4",
X"FD8F",
X"F92A",
X"F4C5",
X"F060",
X"EC78",
X"E890",
X"E525",
X"E1BA",
X"DECC",
X"DBDE",
X"D9EA",
X"D7F6",
X"D67F",
X"D585",
X"D508",
X"D585",
X"D602",
X"D6FC",
X"D873",
X"D9EA",
X"DC5B",
X"DF49",
X"E237",
X"E5A2",
X"E98A",
X"ED72",
X"F1D7",
X"F5BF",
X"FAA1",
X"FF06",
X"036B",
X"07D0",
X"0C35",
X"109A",
X"1482",
X"186A",
X"1C52",
X"1F40",
X"222E",
X"249F",
X"2710",
X"2887",
X"2981",
X"2A7B",
X"2A7B",
X"2A7B",
X"2981",
X"280A",
X"2693",
X"249F",
X"21B1",
X"1EC3",
X"1B58",
X"17ED",
X"1405",
X"0FA0",
X"0B3B",
X"06D6",
X"0271",
X"FD8F",
X"F92A",
X"F4C5",
X"F060",
X"EBFB",
X"E813",
X"E42B",
X"E0C0",
X"DDD2",
X"DB61",
X"D8F0",
X"D6FC",
X"D602",
X"D508",
X"D48B",
X"D508",
X"D585",
X"D67F",
X"D873",
X"DA67",
X"DCD8",
X"DFC6",
X"E331",
X"E719",
X"EB01",
X"EEE9",
X"F34E",
X"F830",
X"FC95",
X"0177",
X"05DC",
X"0ABE",
X"0F23",
X"1388",
X"1770",
X"1B58",
X"1EC3",
X"21B1",
X"249F",
X"2693",
X"2887",
X"29FE",
X"2AF8",
X"2AF8",
X"2AF8",
X"29FE",
X"2904",
X"278D",
X"251C",
X"22AB",
X"1FBD",
X"1C52",
X"186A",
X"1482",
X"101D",
X"0BB8",
X"06D6",
X"0271",
X"FD8F",
X"F8AD",
X"F448",
X"EF66",
X"EB7E",
X"E719",
X"E331",
X"DFC6",
X"DCD8",
X"DA67",
X"D7F6",
X"D67F",
X"D508",
X"D48B",
X"D40E",
X"D48B",
X"D585",
X"D67F",
X"D873",
X"DAE4",
X"DDD2",
X"E0C0",
X"E4A8",
X"E890",
X"EC78",
X"F0DD",
X"F5BF",
X"FA24",
X"FF06",
X"03E8",
X"08CA",
X"0DAC",
X"1211",
X"1676",
X"1A5E",
X"1DC9",
X"2134",
X"2422",
X"2693",
X"2887",
X"29FE",
X"2AF8",
X"2B75",
X"2B75",
X"2AF8",
X"2981",
X"280A",
X"2616",
X"2328",
X"203A",
X"1CCF",
X"18E7",
X"1482",
X"101D",
X"0BB8",
X"06D6",
X"01F4",
X"FD12",
X"F830",
X"F34E",
X"EEE9",
X"EA84",
X"E61F",
X"E237",
X"DECC",
X"DBDE",
X"D96D",
X"D6FC",
X"D585",
X"D48B",
X"D391",
X"D391",
X"D40E",
X"D585",
X"D6FC",
X"D8F0",
X"DB61",
X"DECC",
X"E237",
X"E61F",
X"EA07",
X"EE6C",
X"F34E",
X"F830",
X"FD12",
X"01F4",
X"06D6",
X"0BB8",
X"109A",
X"14FF",
X"1964",
X"1D4C",
X"20B7",
X"23A5",
X"2693",
X"2887",
X"2A7B",
X"2B75",
X"2BF2",
X"2BF2",
X"2B75",
X"2A7B",
X"2887",
X"2693",
X"23A5",
X"20B7",
X"1D4C",
X"1964",
X"14FF",
X"109A",
X"0BB8",
X"06D6",
X"01F4",
X"FC95",
X"F7B3",
X"F2D1",
X"EDEF",
X"E98A",
X"E525",
X"E13D",
X"DDD2",
X"DAE4",
X"D873",
X"D602",
X"D48B",
X"D391",
X"D314",
X"D391",
X"D40E",
X"D585",
X"D6FC",
X"D96D",
X"DC5B",
X"DFC6",
X"E3AE",
X"E796",
X"EBFB",
X"F0DD",
X"F5BF",
X"FAA1",
X"FF83",
X"04E2",
X"09C4",
X"0EA6",
X"1388",
X"17ED",
X"1BD5",
X"1FBD",
X"2328",
X"2616",
X"2887",
X"2A7B",
X"2B75",
X"2C6F",
X"2C6F",
X"2BF2",
X"2AF8",
X"2981",
X"278D",
X"249F",
X"21B1",
X"1DC9",
X"19E1",
X"157C",
X"1117",
X"0C35",
X"06D6",
X"01F4",
X"FC95",
X"F7B3",
X"F254",
X"ED72",
X"E90D",
X"E4A8",
X"E0C0",
X"DD55",
X"D9EA",
X"D779",
X"D585",
X"D40E",
X"D314",
X"D297",
X"D314",
X"D40E",
X"D585",
X"D779",
X"D9EA",
X"DD55",
X"E0C0",
X"E4A8",
X"E90D",
X"EDEF",
X"F2D1",
X"F7B3",
X"FD12",
X"0271",
X"0753",
X"0CB2",
X"1194",
X"15F9",
X"1ADB",
X"1EC3",
X"222E",
X"2599",
X"280A",
X"2A7B",
X"2BF2",
X"2CEC",
X"2CEC",
X"2CEC",
X"2BF2",
X"2A7B",
X"280A",
X"2599",
X"22AB",
X"1EC3",
X"1ADB",
X"1676",
X"1194",
X"0CB2",
X"0753",
X"01F4",
X"FD12",
X"F7B3",
X"F254",
X"ED72",
X"E890",
X"E42B",
X"E043",
X"DC5B",
X"D96D",
X"D6FC",
X"D48B",
X"D314",
X"D297",
X"D21A",
X"D297",
X"D391",
X"D585",
X"D779",
X"DA67",
X"DDD2",
X"E1BA",
X"E5A2",
X"EA84",
X"EF66",
X"F448",
X"F9A7",
X"FF06",
X"0465",
X"09C4",
X"0F23",
X"1405",
X"186A",
X"1CCF",
X"20B7",
X"249F",
X"278D",
X"29FE",
X"2B75",
X"2CEC",
X"2D69",
X"2D69",
X"2CEC",
X"2B75",
X"2981",
X"2710",
X"23A5",
X"203A",
X"1C52",
X"17ED",
X"130B",
X"0DAC",
X"084D",
X"02EE",
X"FD8F",
X"F830",
X"F2D1",
X"EDEF",
X"E90D",
X"E42B",
X"E043",
X"DC5B",
X"D8F0",
X"D67F",
X"D40E",
X"D297",
X"D21A",
X"D19D",
X"D21A",
X"D391",
X"D508",
X"D779",
X"DA67",
X"DDD2",
X"E1BA",
X"E61F",
X"EB01",
X"F060",
X"F542",
X"FB1E",
X"007D",
X"05DC",
X"0B3B",
X"109A",
X"15F9",
X"1A5E",
X"1EC3",
X"22AB",
X"2616",
X"2904",
X"2AF8",
X"2CEC",
X"2DE6",
X"2DE6",
X"2D69",
X"2C6F",
X"2AF8",
X"2887",
X"2599",
X"222E",
X"1E46",
X"19E1",
X"14FF",
X"0FA0",
X"0A41",
X"04E2",
X"FF83",
X"F9A7",
X"F448",
X"EEE9",
X"E98A",
X"E525",
X"E0C0",
X"DCD8",
X"D96D",
X"D67F",
X"D40E",
X"D297",
X"D19D",
X"D120",
X"D19D",
X"D314",
X"D48B",
X"D6FC",
X"D9EA",
X"DDD2",
X"E1BA",
X"E61F",
X"EB01",
X"F060",
X"F5BF",
X"FB9B",
X"00FA",
X"06D6",
X"0C35",
X"1194",
X"16F3",
X"1BD5",
X"203A",
X"2422",
X"2710",
X"29FE",
X"2BF2",
X"2D69",
X"2E63",
X"2E63",
X"2DE6",
X"2C6F",
X"2A7B",
X"280A",
X"249F",
X"20B7",
X"1C52",
X"17ED",
X"128E",
X"0D2F",
X"07D0",
X"01F4",
X"FC18",
X"F63C",
X"F0DD",
X"EB7E",
X"E69C",
X"E1BA",
X"DDD2",
X"D9EA",
X"D6FC",
X"D40E",
X"D297",
X"D120",
X"D0A3",
X"D120",
X"D21A",
X"D391",
X"D602",
X"D8F0",
X"DCD8",
X"E0C0",
X"E5A2",
X"EA84",
X"EFE3",
X"F542",
X"FB1E",
X"00FA",
X"06D6",
X"0C35",
X"1211",
X"16F3",
X"1BD5",
X"20B7",
X"249F",
X"280A",
X"2A7B",
X"2CEC",
X"2DE6",
X"2EE0",
X"2EE0",
X"2DE6",
X"2C6F",
X"2A7B",
X"278D",
X"2422",
X"203A",
X"1B58",
X"1676",
X"1117",
X"0BB8",
X"05DC",
X"0000",
X"FA24",
X"F448",
X"EE6C",
X"E90D",
X"E42B",
X"DFC6",
X"DB61",
X"D7F6",
X"D508",
X"D314",
X"D120",
X"D0A3",
X"D0A3",
X"D120",
X"D297",
X"D48B",
X"D779",
X"DAE4",
X"DECC",
X"E3AE",
X"E890",
X"EDEF",
X"F3CB",
X"F9A7",
X"FF83",
X"055F",
X"0B3B",
X"1117",
X"1676",
X"1B58",
X"203A",
X"2422",
X"280A",
X"2AF8",
X"2CEC",
X"2E63",
X"2F5D",
X"2F5D",
X"2E63",
X"2CEC",
X"2AF8",
X"280A",
X"2422",
X"203A",
X"1B58",
X"1676",
X"1117",
X"0B3B",
X"055F",
X"FF06",
X"F92A",
X"F34E",
X"ED72",
X"E813",
X"E2B4",
X"DE4F",
X"DA67",
X"D6FC",
X"D40E",
X"D21A",
X"D0A3",
X"D026",
X"D026",
X"D120",
X"D314",
X"D585",
X"D873",
X"DC5B",
X"E0C0",
X"E5A2",
X"EB01",
X"F060",
X"F63C",
X"FC95",
X"0271",
X"08CA",
X"0EA6",
X"1482",
X"19E1",
X"1EC3",
X"2328",
X"2710",
X"29FE",
X"2CEC",
X"2E63",
X"2F5D",
X"2FDA",
X"2F5D",
X"2DE6",
X"2BF2",
X"2904",
X"2599",
X"2134",
X"1CCF",
X"1770",
X"1211",
X"0C35",
X"05DC",
X"FF83",
X"F9A7",
X"F34E",
X"ED72",
X"E813",
X"E2B4",
X"DDD2",
X"D9EA",
X"D67F",
X"D391",
X"D19D",
X"D026",
X"CFA9",
X"CFA9",
X"D0A3",
X"D297",
X"D585",
X"D8F0",
X"DCD8",
X"E13D",
X"E69C",
X"EBFB",
X"F1D7",
X"F7B3",
X"FE0C",
X"0465",
X"0ABE",
X"109A",
X"1676",
X"1BD5",
X"20B7",
X"251C",
X"2887",
X"2B75",
X"2DE6",
X"2F5D",
X"3057",
X"2FDA",
X"2EE0",
X"2D69",
X"2AF8",
X"278D",
X"23A5",
X"1F40",
X"19E1",
X"1482",
X"0EA6",
X"084D",
X"01F4",
X"FB9B",
X"F542",
X"EF66",
X"E98A",
X"E42B",
X"DECC",
X"DA67",
X"D6FC",
X"D391",
X"D19D",
X"CFA9",
X"CF2C",
X"CF2C",
X"D026",
X"D21A",
X"D48B",
X"D7F6",
X"DBDE",
X"E0C0",
X"E5A2",
X"EB7E",
X"F15A",
X"F7B3",
X"FE0C",
X"0465",
X"0ABE",
X"1117",
X"16F3",
X"1C52",
X"2134",
X"2599",
X"2981",
X"2C6F",
X"2EE0",
X"2FDA",
X"30D4",
X"3057",
X"2F5D",
X"2D69",
X"2A7B",
X"2710",
X"22AB",
X"1DC9",
X"186A",
X"128E",
X"0CB2",
X"0659",
X"FF83",
X"F92A",
X"F2D1",
X"EC78",
X"E719",
X"E1BA",
X"DCD8",
X"D873",
X"D508",
X"D21A",
X"D026",
X"CF2C",
X"CEAF",
X"CF2C",
X"D0A3",
X"D314",
X"D602",
X"D9EA",
X"DE4F",
X"E3AE",
X"E90D",
X"EF66",
X"F5BF",
X"FC18",
X"0271",
X"0947",
X"0FA0",
X"157C",
X"1B58",
X"20B7",
X"251C",
X"2904",
X"2C6F",
X"2EE0",
X"3057",
X"30D4",
X"30D4",
X"2FDA",
X"2DE6",
X"2AF8",
X"278D",
X"2328",
X"1E46",
X"18E7",
X"130B",
X"0CB2",
X"05DC",
X"FF83",
X"F8AD",
X"F254",
X"EBFB",
X"E61F",
X"E0C0",
X"DBDE",
X"D779",
X"D40E",
X"D120",
X"CF2C",
X"CE32",
X"CE32",
X"CF2C",
X"D120",
X"D391",
X"D6FC",
X"DAE4",
X"DFC6",
X"E525",
X"EB01",
X"F15A",
X"F830",
X"FE89",
X"055F",
X"0C35",
X"128E",
X"186A",
X"1E46",
X"2328",
X"278D",
X"2B75",
X"2DE6",
X"3057",
X"3151",
X"3151",
X"30D4",
X"2EE0",
X"2C6F",
X"2904",
X"251C",
X"203A",
X"1ADB",
X"14FF",
X"0EA6",
X"07D0",
X"00FA",
X"FAA1",
X"F3CB",
X"ED72",
X"E719",
X"E13D",
X"DC5B",
X"D7F6",
X"D40E",
X"D120",
X"CF2C",
X"CE32",
X"CDB5",
X"CEAF",
X"D026",
X"D314",
X"D67F",
X"DA67",
X"DF49",
X"E525",
X"EB01",
X"F15A",
X"F830",
X"FF06",
X"05DC",
X"0CB2",
X"130B",
X"1964",
X"1F40",
X"2422",
X"2887",
X"2BF2",
X"2EE0",
X"30D4",
X"31CE",
X"31CE",
X"30D4",
X"2EE0",
X"2BF2",
X"2887",
X"2422",
X"1EC3",
X"1964",
X"130B",
X"0C35",
X"055F",
X"FE89",
X"F7B3",
X"F0DD",
X"EA84",
X"E42B",
X"DECC",
X"D9EA",
X"D585",
X"D21A",
X"CFA9",
X"CE32",
X"CD38",
X"CDB5",
X"CF2C",
X"D19D",
X"D48B",
X"D873",
X"DD55",
X"E2B4",
X"E890",
X"EF66",
X"F63C",
X"FD12",
X"03E8",
X"0ABE",
X"1194",
X"17ED",
X"1E46",
X"2328",
X"280A",
X"2BF2",
X"2EE0",
X"30D4",
X"324B",
X"324B",
X"3151",
X"2F5D",
X"2CEC",
X"2904",
X"249F",
X"1F40",
X"1964",
X"130B",
X"0C35",
X"055F",
X"FE89",
X"F736",
X"F060",
X"E98A",
X"E3AE",
X"DDD2",
X"D8F0",
X"D48B",
X"D19D",
X"CF2C",
X"CDB5",
X"CD38",
X"CDB5",
X"CF2C",
X"D19D",
X"D508",
X"D96D",
X"DE4F",
X"E42B",
X"EA84",
X"F15A",
X"F830",
X"FF83",
X"0659",
X"0DAC",
X"1482",
X"1ADB",
X"20B7",
X"2599",
X"29FE",
X"2DE6",
X"3057",
X"31CE",
X"32C8",
X"324B",
X"30D4",
X"2E63",
X"2AF8",
X"2710",
X"21B1",
X"1C52",
X"15F9",
X"0F23",
X"084D",
X"00FA",
X"F9A7",
X"F254",
X"EB7E",
X"E525",
X"DF49",
X"D9EA",
X"D585",
X"D19D",
X"CF2C",
X"CD38",
X"CCBB",
X"CD38",
X"CE32",
X"D0A3",
X"D40E",
X"D873",
X"DD55",
X"E331",
X"E98A",
X"F060",
X"F7B3",
X"FF06",
X"0659",
X"0DAC",
X"1482",
X"1ADB",
X"20B7",
X"2616",
X"2A7B",
X"2E63",
X"30D4",
X"324B",
X"3345",
X"32C8",
X"30D4",
X"2E63",
X"2AF8",
X"2693",
X"2134",
X"1B58",
X"1482",
X"0DAC",
X"0659",
X"FF06",
X"F7B3",
X"F060",
X"E98A",
X"E331",
X"DD55",
X"D7F6",
X"D391",
X"D026",
X"CDB5",
X"CCBB",
X"CC3E",
X"CD38",
X"CF2C",
X"D21A",
X"D585",
X"DA67",
X"E043",
X"E61F",
X"ECF5",
X"F448",
X"FB9B",
X"02EE",
X"0ABE",
X"1194",
X"186A",
X"1EC3",
X"249F",
X"2981",
X"2D69",
X"3057",
X"324B",
X"3345",
X"3345",
X"31CE",
X"2F5D",
X"2C6F",
X"280A",
X"22AB",
X"1CCF",
X"1676",
X"0F23",
X"07D0",
X"007D",
X"F8AD",
X"F15A",
X"EA07",
X"E3AE",
X"DD55",
X"D7F6",
X"D391",
X"D026",
X"CDB5",
X"CC3E",
X"CBC1",
X"CCBB",
X"CEAF",
X"D19D",
X"D585",
X"DA67",
X"E043",
X"E69C",
X"ED72",
X"F4C5",
X"FC95",
X"03E8",
X"0BB8",
X"130B",
X"19E1",
X"203A",
X"2616",
X"2A7B",
X"2E63",
X"3151",
X"3345",
X"33C2",
X"3345",
X"31CE",
X"2EE0",
X"2B75",
X"2693",
X"2134",
X"1ADB",
X"1405",
X"0C35",
X"04E2",
X"FD12",
X"F542",
X"EDEF",
X"E719",
X"E043",
X"DA67",
X"D585",
X"D19D",
X"CE32",
X"CC3E",
X"CBC1",
X"CBC1",
X"CD38",
X"D026",
X"D391",
X"D873",
X"DDD2",
X"E42B",
X"EB01",
X"F254",
X"FA24",
X"01F4",
X"09C4",
X"1117",
X"186A",
X"1EC3",
X"249F",
X"29FE",
X"2DE6",
X"3151",
X"3345",
X"343F",
X"33C2",
X"324B",
X"2FDA",
X"2BF2",
X"278D",
X"21B1",
X"1B58",
X"1482",
X"0D2F",
X"055F",
X"FD12",
X"F542",
X"EDEF",
X"E69C",
X"DFC6",
X"D9EA",
X"D508",
X"D0A3",
X"CDB5",
X"CBC1",
X"CB44",
X"CBC1",
X"CD38",
X"D026",
X"D40E",
X"D8F0",
X"DECC",
X"E525",
X"EC78",
X"F3CB",
X"FB9B",
X"03E8",
X"0BB8",
X"130B",
X"1A5E",
X"2134",
X"2710",
X"2BF2",
X"2FDA",
X"324B",
X"343F",
X"34BC",
X"33C2",
X"31CE",
X"2EE0",
X"2A7B",
X"251C",
X"1F40",
X"186A",
X"1117",
X"0947",
X"00FA",
X"F92A",
X"F15A",
X"E98A",
X"E2B4",
X"DC5B",
X"D67F",
X"D21A",
X"CEAF",
X"CC3E",
X"CAC7",
X"CAC7",
X"CC3E",
X"CEAF",
X"D21A",
X"D6FC",
X"DCD8",
X"E331",
X"EA07",
X"F1D7",
X"FA24",
X"01F4",
X"0A41",
X"1211",
X"1964",
X"203A",
X"2616",
X"2B75",
X"2F5D",
X"32C8",
X"343F",
X"34BC",
X"343F",
X"324B",
X"2F5D",
X"2AF8",
X"2599",
X"1F40",
X"186A",
X"1117",
X"0947",
X"00FA",
X"F8AD",
X"F0DD",
X"E90D",
X"E1BA",
X"DB61",
X"D602",
X"D120",
X"CDB5",
X"CB44",
X"CA4A",
X"CAC7",
X"CC3E",
X"CF2C",
X"D314",
X"D7F6",
X"DDD2",
X"E4A8",
X"EBFB",
X"F448",
X"FC18",
X"0465",
X"0CB2",
X"1482",
X"1BD5",
X"22AB",
X"2887",
X"2D69",
X"3151",
X"33C2",
X"3539",
X"3539",
X"33C2",
X"3151",
X"2D69",
X"2887",
X"22AB",
X"1C52",
X"14FF",
X"0CB2",
X"0465",
X"FC18",
X"F3CB",
X"EBFB",
X"E42B",
X"DD55",
X"D779",
X"D297",
X"CEAF",
X"CBC1",
X"CA4A",
X"CA4A",
X"CB44",
X"CDB5",
X"D19D",
X"D67F",
X"DC5B",
X"E2B4",
X"EA84",
X"F254",
X"FAA1",
X"02EE",
X"0B3B",
X"1388",
X"1B58",
X"222E",
X"280A",
X"2D69",
X"3151",
X"33C2",
X"3539",
X"35B6",
X"343F",
X"31CE",
X"2DE6",
X"2904",
X"2328",
X"1C52",
X"1482",
X"0CB2",
X"0465",
X"FB9B",
X"F34E",
X"EB01",
X"E3AE",
X"DC5B",
X"D67F",
X"D19D",
X"CDB5",
X"CB44",
X"C9CD",
X"C9CD",
X"CB44",
X"CE32",
X"D21A",
X"D779",
X"DD55",
X"E4A8",
X"EC78",
X"F4C5",
X"FD12",
X"05DC",
X"0E29",
X"1676",
X"1DC9",
X"249F",
X"2A7B",
X"2F5D",
X"32C8",
X"3539",
X"3633",
X"35B6",
X"33C2",
X"3057",
X"2BF2",
X"2693",
X"1FBD",
X"186A",
X"109A",
X"084D",
X"FF83",
X"F6B9",
X"EE6C",
X"E69C",
X"DECC",
X"D873",
X"D314",
X"CEAF",
X"CBC1",
X"C9CD",
X"C950",
X"CA4A",
X"CCBB",
X"D0A3",
X"D585",
X"DB61",
X"E2B4",
X"EA84",
X"F2D1",
X"FB1E",
X"03E8",
X"0CB2",
X"14FF",
X"1CCF",
X"23A5",
X"29FE",
X"2EE0",
X"32C8",
X"3539",
X"3633",
X"35B6",
X"343F",
X"30D4",
X"2C6F",
X"2710",
X"203A",
X"18E7",
X"109A",
X"07D0",
X"FF06",
X"F63C",
X"EDEF",
X"E5A2",
X"DE4F",
X"D779",
X"D21A",
X"CDB5",
X"CAC7",
X"C950",
X"C950",
X"CA4A",
X"CD38",
X"D120",
X"D67F",
X"DCD8",
X"E42B",
X"EBFB",
X"F4C5",
X"FD8F",
X"0659",
X"0F23",
X"1770",
X"1F40",
X"2616",
X"2BF2",
X"30D4",
X"343F",
X"3633",
X"36B0",
X"35B6",
X"3345",
X"2F5D",
X"2A7B",
X"2422",
X"1D4C",
X"14FF",
X"0CB2",
X"03E8",
X"FAA1",
X"F1D7",
X"E98A",
X"E13D",
X"DA67",
X"D40E",
X"CF2C",
X"CBC1",
X"C950",
X"C8D3",
X"C950",
X"CBC1",
X"CF2C",
X"D40E",
X"DA67",
X"E13D",
X"E98A",
X"F1D7",
X"FB1E",
X"03E8",
X"0D2F",
X"157C",
X"1DC9",
X"251C",
X"2AF8",
X"3057",
X"33C2",
X"3633",
X"372D",
X"3633",
X"343F",
X"3057",
X"2B75",
X"251C",
X"1E46",
X"15F9",
X"0D2F",
X"0465",
X"FB1E",
X"F1D7",
X"E98A",
X"E13D",
X"D9EA",
X"D40E",
X"CEAF",
X"CB44",
X"C8D3",
X"C856",
X"C950",
X"CBC1",
X"CF2C",
X"D48B",
X"DAE4",
X"E237",
X"EA84",
X"F34E",
X"FC95",
X"05DC",
X"0F23",
X"1770",
X"1FBD",
X"2693",
X"2CEC",
X"31CE",
X"3539",
X"36B0",
X"372D",
X"3633",
X"3345",
X"2F5D",
X"2981",
X"2328",
X"1B58",
X"130B",
X"09C4",
X"007D",
X"F736",
X"EE6C",
X"E5A2",
X"DDD2",
X"D6FC",
X"D120",
X"CCBB",
X"C9CD",
X"C856",
X"C856",
X"C9CD",
X"CD38",
X"D19D",
X"D7F6",
X"DECC",
X"E719",
X"EFE3",
X"F8AD",
X"0271",
X"0BB8",
X"1482",
X"1D4C",
X"249F",
X"2B75",
X"3057",
X"343F",
X"36B0",
X"37AA",
X"36B0",
X"34BC",
X"30D4",
X"2B75",
X"249F",
X"1D4C",
X"1482",
X"0BB8",
X"0271",
X"F8AD",
X"EF66",
X"E69C",
X"DE4F",
X"D779",
X"D120",
X"CCBB",
X"C950",
X"C7D9",
X"C7D9",
X"C950",
X"CCBB",
X"D19D",
X"D779",
X"DECC",
X"E719",
X"EFE3",
X"F92A",
X"02EE",
X"0C35",
X"157C",
X"1DC9",
X"2599",
X"2BF2",
X"3151",
X"3539",
X"372D",
X"3827",
X"36B0",
X"343F",
X"2FDA",
X"2A7B",
X"23A5",
X"1B58",
X"128E",
X"0947",
X"0000",
X"F63C",
X"ECF5",
X"E42B",
X"DBDE",
X"D508",
X"CF2C",
X"CB44",
X"C856",
X"C75C",
X"C7D9",
X"CA4A",
X"CE32",
X"D391",
X"DA67",
X"E1BA",
X"EA84",
X"F3CB",
X"FD8F",
X"0753",
X"1117",
X"19E1",
X"222E",
X"2981",
X"2F5D",
X"33C2",
X"36B0",
X"3827",
X"37AA",
X"35B6",
X"324B",
X"2CEC",
X"2693",
X"1EC3",
X"15F9",
X"0CB2",
X"02EE",
X"F92A",
X"EF66",
X"E61F",
X"DDD2",
X"D67F",
X"D0A3",
X"CBC1",
X"C8D3",
X"C75C",
X"C75C",
X"C950",
X"CD38",
X"D21A",
X"D8F0",
X"E043",
X"E90D",
X"F2D1",
X"FC95",
X"0659",
X"101D",
X"1964",
X"21B1",
X"2904",
X"2F5D",
X"343F",
X"372D",
X"38A4",
X"3827",
X"3633",
X"324B",
X"2CEC",
X"2693",
X"1EC3",
X"157C",
X"0C35",
X"0271",
X"F830",
X"EE6C",
X"E525",
X"DCD8",
X"D585",
X"CF2C",
X"CAC7",
X"C7D9",
X"C6DF",
X"C75C",
X"C9CD",
X"CDB5",
X"D314",
X"DA67",
X"E237",
X"EB7E",
X"F542",
X"FF06",
X"0947",
X"130B",
X"1C52",
X"249F",
X"2B75",
X"3151",
X"35B6",
X"3827",
X"3921",
X"3827",
X"3539",
X"30D4",
X"2A7B",
X"2328",
X"1ADB",
X"1194",
X"0753",
X"FD8F",
X"F34E",
X"E98A",
X"E0C0",
X"D873",
X"D19D",
X"CC3E",
X"C8D3",
X"C6DF",
X"C662",
X"C856",
X"CBC1",
X"D0A3",
X"D779",
X"DF49",
X"E813",
X"F1D7",
X"FB9B",
X"05DC",
X"101D",
X"19E1",
X"222E",
X"29FE",
X"3057",
X"3539",
X"3827",
X"3921",
X"38A4",
X"3633",
X"31CE",
X"2BF2",
X"251C",
X"1C52",
X"130B",
X"0947",
X"FE89",
X"F448",
X"EA84",
X"E13D",
X"D8F0",
X"D21A",
X"CC3E",
X"C856",
X"C662",
X"C662",
X"C7D9",
X"CB44",
X"D0A3",
X"D6FC",
X"DF49",
X"E813",
X"F1D7",
X"FC95",
X"06D6",
X"1117",
X"1ADB",
X"2328",
X"2AF8",
X"3151",
X"35B6",
X"38A4",
X"399E",
X"38A4",
X"35B6",
X"3151",
X"2AF8",
X"23A5",
X"1ADB",
X"1117",
X"06D6",
X"FC18",
X"F1D7",
X"E796",
X"DECC",
X"D67F",
X"CFA9",
X"CAC7",
X"C75C",
X"C5E5",
X"C662",
X"C856",
X"CCBB",
X"D297",
X"D9EA",
X"E2B4",
X"EBFB",
X"F63C",
X"00FA",
X"0B3B",
X"157C",
X"1EC3",
X"278D",
X"2E63",
X"33C2",
X"37AA",
X"399E",
X"399E",
X"37AA",
X"33C2",
X"2E63",
X"2710",
X"1EC3",
X"14FF",
X"0ABE",
X"0000",
X"F5BF",
X"EB01",
X"E1BA",
X"D8F0",
X"D19D",
X"CBC1",
X"C7D9",
X"C5E5",
X"C5E5",
X"C75C",
X"CB44",
X"D0A3",
X"D7F6",
X"E043",
X"EA07",
X"F448",
X"FE89",
X"0947",
X"1405",
X"1DC9",
X"2693",
X"2DE6",
X"33C2",
X"37AA",
X"399E",
X"3A1B",
X"3827",
X"343F",
X"2EE0",
X"278D",
X"1F40",
X"157C",
X"0B3B",
X"007D",
X"F5BF",
X"EB01",
X"E13D",
X"D873",
X"D120",
X"CB44",
X"C75C",
X"C568",
X"C568",
X"C75C",
X"CB44",
X"D120",
X"D873",
X"E13D",
X"EB01",
X"F5BF",
X"007D",
X"0B3B",
X"15F9",
X"1FBD",
X"280A",
X"2F5D",
X"34BC",
X"38A4",
X"3A98",
X"3A1B",
X"37AA",
X"3345",
X"2D69",
X"2599",
X"1C52",
X"128E",
X"07D0",
X"FC95",
X"F1D7",
X"E719",
X"DDD2",
X"D585",
X"CEAF",
X"C950",
X"C5E5",
X"C4EB",
X"C5E5",
X"C8D3",
X"CDB5",
X"D40E",
X"DC5B",
X"E5A2",
X"F060",
X"FB1E",
X"0659",
X"1117",
X"1B58",
X"249F",
X"2C6F",
X"3345",
X"37AA",
X"3A1B",
X"3A98",
X"3921",
X"3539",
X"2FDA",
X"2887",
X"1FBD",
X"15F9",
X"0B3B",
X"0000",
X"F4C5",
X"EA07",
X"E043",
X"D779",
X"CFA9",
X"CA4A",
X"C662",
X"C4EB",
X"C4EB",
X"C7D9",
X"CC3E",
X"D297",
X"DAE4",
X"E42B",
X"EE6C",
X"F9A7",
X"04E2",
X"101D",
X"1A5E",
X"2422",
X"2C6F",
X"32C8",
X"37AA",
X"3A98",
X"3B15",
X"399E",
X"35B6",
X"3057",
X"2904",
X"1FBD",
X"15F9",
X"0B3B",
X"FF83",
X"F448",
X"E98A",
X"DF49",
X"D67F",
X"CF2C",
X"C950",
X"C5E5",
X"C46E",
X"C4EB",
X"C7D9",
X"CCBB",
X"D391",
X"DBDE",
X"E5A2",
X"F060",
X"FB9B",
X"0753",
X"1211",
X"1CCF",
X"2616",
X"2E63",
X"34BC",
X"38A4",
X"3B15",
X"3B15",
X"3921",
X"34BC",
X"2E63",
X"2616",
X"1CCF",
X"1211",
X"06D6",
X"FB9B",
X"EFE3",
X"E525",
X"DB61",
X"D314",
X"CC3E",
X"C75C",
X"C46E",
X"C3F1",
X"C5E5",
X"C9CD",
X"CFA9",
X"D779",
X"E0C0",
X"EB01",
X"F63C",
X"01F4",
X"0D2F",
X"186A",
X"22AB",
X"2B75",
X"324B",
X"37AA",
X"3A98",
X"3B92",
X"3A1B",
X"36B0",
X"30D4",
X"2981",
X"203A",
X"15F9",
X"0ABE",
X"FF06",
X"F34E",
X"E813",
X"DDD2",
X"D508",
X"CDB5",
X"C856",
X"C4EB",
X"C3F1",
X"C4EB",
X"C856",
X"CE32",
X"D585",
X"DECC",
X"E90D",
X"F448",
X"0000",
X"0BB8",
X"16F3",
X"21B1",
X"2A7B",
X"31CE",
X"37AA",
X"3B15",
X"3C0F",
X"3A98",
X"372D",
X"3151",
X"29FE",
X"20B7",
X"15F9",
X"0ABE",
X"FF06",
X"F2D1",
X"E796",
X"DD55",
X"D40E",
X"CCBB",
X"C75C",
X"C46E",
X"C374",
X"C4EB",
X"C8D3",
X"CEAF",
X"D67F",
X"DFC6",
X"EA84",
X"F63C",
X"0271",
X"0E29",
X"1964",
X"23A5",
X"2C6F",
X"33C2",
X"38A4",
X"3B92",
X"3C0F",
X"3A1B",
X"3633",
X"2FDA",
X"278D",
X"1DC9",
X"128E",
X"06D6",
X"FAA1",
X"EEE9",
X"E3AE",
X"D96D",
X"D120",
X"CA4A",
X"C5E5",
X"C374",
X"C374",
X"C5E5",
X"CAC7",
X"D19D",
X"DA67",
X"E4A8",
X"EFE3",
X"FC18",
X"084D",
X"1405",
X"1EC3",
X"2887",
X"30D4",
X"372D",
X"3B15",
X"3C8C",
X"3B92",
X"3827",
X"32C8",
X"2AF8",
X"21B1",
X"16F3",
X"0B3B",
X"FF06",
X"F2D1",
X"E796",
X"DCD8",
X"D391",
X"CBC1",
X"C662",
X"C374",
X"C2F7",
X"C4EB",
X"C950",
X"CFA9",
X"D7F6",
X"E237",
X"ED72",
X"F9A7",
X"05DC",
X"1194",
X"1D4C",
X"2710",
X"2FDA",
X"3633",
X"3A98",
X"3C8C",
X"3C0F",
X"3921",
X"33C2",
X"2BF2",
X"22AB",
X"17ED",
X"0C35",
X"0000",
X"F34E",
X"E796",
X"DCD8",
X"D391",
X"CBC1",
X"C662",
X"C374",
X"C27A",
X"C46E",
X"C8D3",
X"CFA9",
X"D873",
X"E2B4",
X"EE6C",
X"FAA1",
X"06D6",
X"130B",
X"1EC3",
X"2887",
X"3151",
X"37AA",
X"3B92",
X"3D09",
X"3C0F",
X"38A4",
X"32C8",
X"2A7B",
X"20B7",
X"157C",
X"0947",
X"FC95",
X"F060",
X"E4A8",
X"D9EA",
X"D0A3",
X"C9CD",
X"C4EB",
X"C27A",
X"C2F7",
X"C568",
X"CAC7",
X"D21A",
X"DBDE",
X"E69C",
X"F2D1",
X"FF83",
X"0BB8",
X"17ED",
X"2328",
X"2C6F",
X"343F",
X"399E",
X"3C8C",
X"3D09",
X"3B15",
X"3633",
X"2EE0",
X"2616",
X"1B58",
X"0F23",
X"02EE",
X"F63C",
X"E98A",
X"DE4F",
X"D48B",
X"CC3E",
X"C662",
X"C2F7",
X"C1FD",
X"C3F1",
X"C856",
X"CF2C",
X"D7F6",
X"E2B4",
X"EE6C",
X"FB1E",
X"07D0",
X"1482",
X"203A",
X"2A7B",
X"32C8",
X"38A4",
X"3C8C",
X"3D86",
X"3C0F",
X"37AA",
X"30D4",
X"280A",
X"1DC9",
X"1194",
X"04E2",
X"F830",
X"EB7E",
X"DFC6",
X"D585",
X"CD38",
X"C6DF",
X"C2F7",
X"C1FD",
X"C374",
X"C7D9",
X"CE32",
X"D6FC",
X"E1BA",
X"EDEF",
X"FAA1",
X"07D0",
X"1405",
X"203A",
X"2A7B",
X"32C8",
X"3921",
X"3D09",
X"3E03",
X"3C0F",
X"37AA",
X"30D4",
X"278D",
X"1CCF",
X"109A",
X"03E8",
X"F6B9",
X"EA07",
X"DE4F",
X"D40E",
X"CBC1",
X"C5E5",
X"C27A",
X"C180",
X"C3F1",
X"C856",
X"CFA9",
X"D8F0",
X"E42B",
X"F060",
X"FD8F",
X"0ABE",
X"1770",
X"2328",
X"2CEC",
X"3539",
X"3A98",
X"3D86",
X"3E03",
X"3B15",
X"35B6",
X"2DE6",
X"2422",
X"18E7",
X"0C35",
X"FF06",
X"F1D7",
X"E525",
X"D9EA",
X"D026",
X"C8D3",
X"C374",
X"C180",
X"C1FD"


 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= Jump_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;