library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity yacht_150_30-2_object is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end yacht_150_30-2_object;

architecture behav of yacht_150_30-2_object is

constant object_X_size : integer := 150;
constant object_Y_size : integer := 30;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"00", x"00", x"00", x"00", x"24", x"6D", x"92", x"B6", x"B6", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"49", x"69", x"49", x"49", x"49", x"49", x"49", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"FF", x"FF", x"DB", x"B6", x"92", x"6D", x"6D", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"24", x"D1", x"00", x"24", x"6D", x"6D", x"92", x"92", x"6D", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"D6", x"D6", x"D6", x"D6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"D7", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"8D", x"6D", x"6D", x"49", x"49", x"49", x"24", x"00", x"00", x"FF", x"DB", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"20", x"69", x"8D", x"8D", x"D6", x"DB", x"FB", x"DB", x"B6", x"B6", x"D7", x"D7", x"D6", x"D6", x"D6", x"D6", x"D6", x"B6", x"B6", x"B6", x"B6", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B2", x"B6", x"D6", x"B6", x"D6", x"D6", x"D6", x"DA", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"B6", x"B6", x"B6", x"92", x"6D", x"6D", x"24", x"00", x"00", x"FF", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"68", x"B1", x"D1", x"B1", x"B2", x"D6", x"B6", x"B6", x"B6", x"B6", x"B2", x"B2", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"DB", x"DB", x"FB", x"FF", x"FF", x"FB", x"DB", x"DB", x"DB", x"B6", x"92", x"8D", x"49", x"00", x"00", x"FF", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"24", x"8D", x"B1", x"B1", x"B1", x"B1", x"AD", x"B1", x"B1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"D6", x"DA", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"D6", x"B6", x"B6", x"B6", x"B2", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B2", x"B2", x"B6", x"B6", x"B6", x"D6", x"D6", x"DA", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"D6", x"B6", x"B6", x"B6", x"D6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"DA", x"DA", x"DA", x"DA", x"DA", x"DA", x"DA", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D5", x"D5", x"D1", x"D1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D6", x"D6", x"DA", x"DB", x"FB", x"FF", x"FF", x"FB", x"DB", x"DB", x"B6", x"92", x"8D", x"49", x"00", x"FF", x"B6", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"48", x"B1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B2", x"D1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"D7", x"D7", x"DB", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"FB", x"FF", x"DB", x"92", x"92", x"92", x"72", x"6E", x"6E", x"4D", x"4D", x"4D", x"49", x"49", x"49", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"DA", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D5", x"D1", x"B1", x"B1", x"D1", x"D1", x"D6", x"D6", x"DA", x"FB", x"FF", x"FF", x"FB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"FF", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"68", x"B1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B2", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"FF", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"FF", x"DB", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"25", x"01", x"25", x"25", x"29", x"29", x"29", x"29", x"49", x"49", x"49", x"49", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DA", x"D6", x"DA", x"DB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DB", x"DB", x"FB", x"FB", x"FF", x"FF", x"FB", x"FA", x"D6", x"D1", x"B1", x"D1", x"B1", x"B1", x"B1", x"D1", x"D6", x"D6", x"DA", x"FB", x"FF", x"FF", x"DB", x"DB", x"B6", x"6D", x"24", x"00", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"69", x"D1", x"D1", x"D1", x"B1", x"B1", x"B2", x"D6", x"D6", x"B6", x"B2", x"B2", x"B1", x"B1", x"D6", x"DB", x"D7", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6E", x"25", x"25", x"25", x"49", x"49", x"49", x"49", x"49", x"49", x"4E", x"4E", x"49", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"DB", x"DB", x"DB", x"DA", x"DA", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"DA", x"DB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B2", x"D6", x"DA", x"FB", x"FF", x"FB", x"DB", x"B6", x"92", x"49", x"00", x"D6", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"8D", x"D1", x"D1", x"D1", x"B1", x"B6", x"B6", x"DB", x"DB", x"D6", x"B6", x"B6", x"B6", x"B1", x"D6", x"FF", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"49", x"29", x"25", x"49", x"4D", x"6D", x"6D", x"4D", x"4D", x"6D", x"6E", x"6E", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FB", x"FB", x"DB", x"DB", x"DA", x"DA", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"D6", x"FB", x"FF", x"FF", x"DB", x"B6", x"92", x"49", x"00", x"B6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"8D", x"D1", x"D1", x"B1", x"B2", x"B6", x"D6", x"FA", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"25", x"25", x"49", x"6D", x"72", x"72", x"6E", x"6D", x"6D", x"6D", x"72", x"92", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"D1", x"D6", x"DB", x"FF", x"FF", x"DB", x"B6", x"92", x"00", x"DB", x"49", x"00", x"00", x"00", x"00", x"00"),
(x"8D", x"B1", x"B1", x"B1", x"B6", x"B7", x"D6", x"FB", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"25", x"25", x"24", x"24", x"49", x"92", x"92", x"92", x"6E", x"6D", x"6D", x"6E", x"72", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"FB", x"FF", x"FB", x"D6", x"92", x"24", x"FF", x"49", x"00", x"00", x"00"),
(x"8D", x"D1", x"D1", x"D1", x"B6", x"B6", x"DA", x"FB", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"24", x"24", x"24", x"24", x"49", x"92", x"B6", x"92", x"72", x"6D", x"6D", x"6E", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"D1", x"D6", x"DA", x"FF", x"FF", x"DB", x"92", x"24", x"DB", x"49", x"00"),
(x"8D", x"D1", x"D1", x"D1", x"B6", x"B6", x"DA", x"FA", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"24", x"24", x"49", x"6D", x"92", x"96", x"92", x"6D", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"D1", x"DA", x"FF", x"FF", x"DB", x"92", x"24", x"92"),
(x"8D", x"D1", x"D1", x"D1", x"B6", x"B6", x"DA", x"FA", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"92", x"96", x"92", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"DA", x"FF", x"FF", x"D7", x"6D"),
(x"8D", x"D1", x"B1", x"B1", x"B6", x"B6", x"FA", x"FA", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"6D", x"6D", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"24", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D6", x"FF", x"FF", x"B6"),
(x"8D", x"D1", x"D1", x"D1", x"B6", x"B6", x"FA", x"FB", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"29", x"49", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"24", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"FB", x"FF", x"B6"),
(x"8D", x"D1", x"D1", x"B1", x"B6", x"B6", x"FA", x"FA", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"49", x"6D", x"92", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"8E", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"D1", x"D1", x"D1", x"D1", x"B1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"FB", x"FF", x"DB", x"92"),
(x"8D", x"B1", x"B1", x"B1", x"B6", x"B6", x"FA", x"FA", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"49", x"6D", x"6D", x"6E", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"DA", x"FF", x"FB", x"B6", x"92", x"00"),
(x"8D", x"D1", x"D1", x"B1", x"B6", x"B6", x"DA", x"FA", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"24", x"49", x"4D", x"4D", x"6D", x"6D", x"6E", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"DB", x"FF", x"FB", x"D6", x"92", x"00", x"B6", x"24"),
(x"8D", x"D1", x"D1", x"D1", x"B2", x"B6", x"DA", x"FB", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"24", x"49", x"4D", x"4D", x"4D", x"6D", x"6D", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"B1", x"B1", x"B1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D6", x"FB", x"FF", x"DB", x"B6", x"92", x"00", x"B6", x"00", x"00", x"00"),
(x"8D", x"D1", x"D1", x"D1", x"B2", x"B6", x"D6", x"FB", x"D6", x"D6", x"D6", x"D6", x"B1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"49", x"49", x"4D", x"4D", x"4D", x"6D", x"4D", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"B1", x"D1", x"D6", x"DB", x"FF", x"FF", x"DB", x"B6", x"6D", x"00", x"B6", x"24", x"00", x"00", x"00", x"00"),
(x"8D", x"D1", x"D1", x"D1", x"B2", x"B6", x"D6", x"FB", x"DA", x"D6", x"D6", x"D6", x"B2", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"4D", x"4D", x"4D", x"72", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D1", x"D6", x"DB", x"FF", x"FF", x"DB", x"B6", x"92", x"6D", x"00", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"8D", x"D1", x"D1", x"D1", x"B1", x"B6", x"B6", x"DB", x"DB", x"D6", x"B6", x"B6", x"B2", x"B1", x"D6", x"FF", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"4D", x"4D", x"4D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"DB", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"DA", x"DA", x"DA", x"DB", x"FF", x"FF", x"FF", x"FF", x"FA", x"D6", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"D6", x"FB", x"FF", x"FF", x"DB", x"B6", x"92", x"6D", x"00", x"FF", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"68", x"B1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B2", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"DB", x"D7", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"25", x"00", x"00", x"24", x"49", x"49", x"49", x"29", x"29", x"49", x"4D", x"4D", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"DA", x"DA", x"DA", x"DB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D6", x"D1", x"D1", x"D1", x"D1", x"D1", x"B1", x"B1", x"D1", x"D6", x"D6", x"DB", x"FF", x"FF", x"FB", x"DB", x"B6", x"92", x"49", x"00", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"68", x"B1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B2", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D5", x"FF", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"FF", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"25", x"29", x"49", x"49", x"49", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"DA", x"DA", x"DA", x"DA", x"D6", x"D6", x"D1", x"D1", x"B1", x"B1", x"D1", x"D1", x"D6", x"D6", x"DA", x"FB", x"FF", x"FF", x"FB", x"DB", x"B6", x"92", x"6D", x"24", x"00", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"24", x"AD", x"D1", x"D1", x"B1", x"B1", x"B1", x"B2", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DB", x"DB", x"DB", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B2", x"B6", x"B6", x"B6", x"D7", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"D7", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"B6", x"FB", x"FB", x"FB", x"FB", x"FB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D5", x"D1", x"D1", x"D1", x"B1", x"B1", x"D1", x"B1", x"D2", x"D6", x"D6", x"DA", x"FB", x"FF", x"FF", x"FB", x"DB", x"DB", x"B6", x"92", x"6D", x"49", x"00", x"FF", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"69", x"B1", x"D1", x"B1", x"B1", x"B1", x"B2", x"B2", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B2", x"B2", x"B2", x"B2", x"B2", x"D6", x"B6", x"B6", x"B6", x"B2", x"B6", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B6", x"B6", x"B6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D5", x"D6", x"D5", x"D1", x"D1", x"D1", x"B1", x"D1", x"D1", x"D1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"D6", x"D6", x"D6", x"DB", x"FB", x"FB", x"FF", x"FF", x"FB", x"DB", x"DB", x"B6", x"92", x"8D", x"49", x"00", x"00", x"FF", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"44", x"8D", x"AD", x"B1", x"D6", x"FF", x"FB", x"DB", x"B6", x"D6", x"D6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B2", x"B2", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"AD", x"AD", x"AD", x"AD", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B2", x"B6", x"D6", x"D6", x"D6", x"D6", x"DA", x"DB", x"DB", x"DB", x"DB", x"FB", x"FB", x"DB", x"DB", x"DB", x"DB", x"B6", x"B6", x"B6", x"92", x"6D", x"49", x"00", x"00", x"FF", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"68", x"00", x"48", x"69", x"92", x"B6", x"B6", x"B6", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B6", x"B6", x"B6", x"B6", x"B6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"DA", x"DA", x"DA", x"D6", x"D6", x"DA", x"DA", x"DA", x"DA", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"D7", x"B6", x"B6", x"B6", x"B6", x"B2", x"92", x"92", x"92", x"6D", x"6D", x"49", x"24", x"00", x"00", x"FF", x"D6", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
(x"00", x"00", x"24", x"48", x"8D", x"FF", x"FF", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"49", x"49", x"49", x"49", x"69", x"6D", x"6D", x"6D", x"6D", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B2", x"B2", x"B2", x"B2", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"8E", x"6D", x"6D", x"6D", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"FF", x"FF", x"DB", x"B2", x"6D", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;
  end process;
end behav;		

--generated with PNGtoVHDL tool by Ben Wellingstein
