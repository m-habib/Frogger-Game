library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity speedboat_150_30_object is
port 	(
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end speedboat_150_30_object;

architecture behav of speedboat_150_30_object is

constant object_X_size : integer := 150;
constant object_Y_size : integer := 30;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"48", x"48", x"48", x"49", x"48", x"48", x"6D", x"6D", x"6C", x"6D", x"6D", x"6C", x"6D", x"6D", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6C", x"44", x"92", x"48", x"44", x"00", x"00"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"24", x"24", x"49", x"49", x"25", x"25", x"25", x"29", x"29", x"49", x"4D", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"8D", x"49", x"48", x"48", x"48", x"48", x"49", x"48", x"49", x"48", x"69", x"48", x"69", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"8D", x"68", x"48", x"FF", x"48", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"2E", x"4E", x"4E", x"92", x"B6", x"DB", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"B6", x"92", x"92", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"92", x"92", x"B6", x"92", x"92", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"B6", x"B6", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"8D", x"68", x"6C", x"68", x"6C", x"68", x"68", x"68", x"68", x"6C", x"6D", x"6D", x"48", x"24"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"29", x"29", x"29", x"2E", x"4E", x"4E", x"6E", x"92", x"B6", x"DB", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"92", x"B6", x"92", x"92", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"B6", x"92", x"92", x"92", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"B6", x"B6", x"B6", x"92", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"91", x"B1", x"B1", x"B1", x"B1", x"B1", x"91", x"8D", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"B6", x"B1", x"B1", x"91", x"91", x"91", x"91", x"91", x"91", x"8D", x"8D", x"8D", x"B1", x"B2", x"92", x"6D", x"48", x"68", x"68", x"6D", x"48", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"96", x"DB", x"DB", x"B6", x"92", x"92", x"B6", x"DB", x"B6", x"B6", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"6D", x"6D", x"92", x"92", x"B6", x"92", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"B2", x"B6", x"B6", x"D6", x"B6", x"D6", x"92", x"49", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"B6", x"8D", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"8C", x"8D", x"92", x"6D", x"68", x"68", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"B6", x"DB", x"DB", x"B6", x"92", x"B6", x"92", x"92", x"92", x"6D", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"24", x"49", x"6D", x"6D", x"6D", x"49", x"49", x"6D", x"6D", x"92", x"6D", x"92", x"92", x"92", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"6D", x"6D", x"6D", x"91", x"92", x"B6", x"B6", x"92", x"92", x"91", x"92", x"91", x"8D", x"6D", x"8D", x"6D", x"91", x"6D", x"6D", x"68", x"68", x"68", x"68", x"68", x"88", x"B2", x"92", x"49", x"68", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"72", x"B6", x"DB", x"DB", x"B6", x"92", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"B6", x"6D", x"24", x"00", x"24", x"24", x"49", x"24", x"24", x"49", x"92", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"6D", x"49", x"2A", x"2A", x"2A", x"4E", x"4E", x"4E", x"4E", x"4E", x"4E", x"4A", x"6E", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"92", x"92", x"92", x"B2", x"B2", x"B2", x"B2", x"92", x"92", x"92", x"92", x"B2", x"B2", x"92", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"92", x"91", x"6D", x"92", x"91", x"68", x"68", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"92", x"B6", x"DB", x"B6", x"B6", x"92", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"6D", x"92", x"49", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"29", x"2A", x"2E", x"4F", x"4F", x"2F", x"4F", x"4F", x"73", x"73", x"73", x"6E", x"6D", x"6C", x"8C", x"6C", x"6C", x"8C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"68", x"6C", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"6C", x"68", x"6D", x"92", x"92", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"29", x"29", x"29", x"2E", x"4E", x"4E", x"6E", x"92", x"B6", x"DB", x"B6", x"92", x"92", x"6D", x"92", x"92", x"92", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"49", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"4E", x"73", x"72", x"8D", x"88", x"88", x"88", x"68", x"88", x"68", x"68", x"44", x"44", x"44", x"44", x"44", x"44", x"68", x"92", x"D6", x"D6", x"B6", x"92", x"91", x"91", x"91", x"91", x"91", x"91", x"B2", x"B6", x"92", x"6D", x"91", x"92", x"B2", x"B2", x"B6", x"B6", x"B6", x"B6", x"88", x"68", x"68", x"8D", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"49", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"96", x"DB", x"DB", x"B6", x"92", x"92", x"B6", x"DB", x"B6", x"B6", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"2F", x"2E", x"2F", x"2F", x"4F", x"73", x"B6", x"AC", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"44", x"44", x"68", x"88", x"8D", x"D6", x"DB", x"B6", x"B6", x"8D", x"48", x"44", x"44", x"44", x"44", x"44", x"48", x"92", x"B6", x"49", x"6E", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"8C", x"68", x"68", x"B6", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"B7", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"B6", x"DB", x"DB", x"B6", x"92", x"92", x"92", x"92", x"92", x"6D", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"2F", x"2F", x"2E", x"2F", x"4F", x"73", x"B6", x"D1", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"8C", x"B6", x"DB", x"B6", x"92", x"92", x"6D", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"92", x"B6", x"49", x"6D", x"92", x"92", x"B6", x"B6", x"B6", x"DB", x"DB", x"DB", x"8C", x"68", x"68", x"B6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"88", x"68", x"68", x"6D", x"91", x"B6", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"92", x"DB", x"DB", x"DB", x"B6", x"92", x"92", x"DB", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"91", x"8D", x"B1", x"B1", x"B1", x"B1", x"B1", x"B1", x"91", x"91", x"B1", x"91", x"D6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"2F", x"2F", x"2F", x"2F", x"4F", x"B6", x"B1", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"88", x"B6", x"DB", x"B6", x"92", x"92", x"6D", x"24", x"24", x"24", x"24", x"24", x"25", x"49", x"92", x"DB", x"92", x"72", x"92", x"92", x"B6", x"DB", x"DB", x"B6", x"B6", x"DB", x"8C", x"88", x"68", x"8C", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"24", x"49", x"49", x"6D", x"49", x"25", x"25", x"29", x"4E", x"4E", x"4E", x"4D", x"92", x"DB", x"DB", x"DB", x"92", x"6D", x"92", x"92", x"92", x"6D", x"B6", x"DB", x"DB", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"68", x"AC", x"8C", x"88", x"88", x"8C", x"88", x"88", x"88", x"8C", x"88", x"B6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"2F", x"2F", x"2E", x"2E", x"4F", x"96", x"8C", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"68", x"B6", x"DB", x"B6", x"B6", x"6D", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"29", x"92", x"B7", x"6E", x"6E", x"6D", x"92", x"DB", x"DB", x"DB", x"8D", x"91", x"DB", x"8C", x"88", x"68", x"8C", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"88", x"68", x"48", x"6D", x"91", x"B6", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"25", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"92", x"DB", x"DB", x"DB", x"B6", x"6D", x"B6", x"DB", x"DB", x"92", x"B6", x"DB", x"DB", x"DB", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"68", x"AC", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8C", x"88", x"B6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"2F", x"4F", x"4E", x"2E", x"2E", x"4E", x"92", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"68", x"B6", x"DB", x"B6", x"B6", x"6D", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"29", x"92", x"B7", x"4E", x"6E", x"92", x"92", x"92", x"B6", x"B6", x"8D", x"91", x"DB", x"8C", x"8C", x"68", x"B6", x"DA", x"DA", x"D6", x"D6", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"24", x"24", x"49", x"49", x"4D", x"25", x"25", x"29", x"4E", x"4E", x"4E", x"4E", x"72", x"DB", x"DB", x"DB", x"B6", x"6D", x"92", x"92", x"92", x"6D", x"B6", x"DB", x"DB", x"DB", x"DB", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"68", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"B6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"4E", x"2E", x"2E", x"4E", x"92", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"68", x"B6", x"DB", x"B6", x"B6", x"6D", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"29", x"92", x"B6", x"49", x"6E", x"6D", x"49", x"92", x"DB", x"DB", x"B6", x"B6", x"DB", x"8D", x"DA", x"B1", x"D6", x"DB", x"DA", x"DA", x"DB", x"DB", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"88", x"68", x"68", x"6D", x"91", x"B6", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"24", x"24", x"49", x"49", x"4D", x"25", x"25", x"29", x"4E", x"4E", x"4E", x"4E", x"72", x"DB", x"DB", x"DB", x"B6", x"6D", x"92", x"92", x"92", x"6D", x"B6", x"DB", x"DB", x"DB", x"DB", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"68", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"B6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"2E", x"4E", x"92", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"68", x"B6", x"DB", x"B6", x"B6", x"6D", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"29", x"92", x"B6", x"49", x"6E", x"6D", x"49", x"92", x"DB", x"DB", x"B6", x"B6", x"DB", x"8D", x"DA", x"B1", x"B1", x"DA", x"B6", x"91", x"B6", x"DA", x"B1", x"91", x"91", x"91", x"B1", x"B1", x"88", x"68", x"68", x"6D", x"91", x"B6", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"25", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"92", x"DB", x"DB", x"DB", x"B6", x"6D", x"B6", x"DB", x"DB", x"92", x"B6", x"DB", x"DB", x"DB", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"68", x"AC", x"8C", x"88", x"8C", x"8C", x"88", x"88", x"88", x"8C", x"88", x"B6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"2E", x"4E", x"92", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"68", x"B6", x"DB", x"B6", x"B6", x"6D", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"29", x"92", x"B7", x"4E", x"6E", x"92", x"6D", x"6D", x"6E", x"B6", x"8D", x"91", x"DB", x"8C", x"8C", x"8C", x"8C", x"8D", x"8C", x"8C", x"8C", x"8D", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"24", x"49", x"49", x"6D", x"49", x"25", x"25", x"29", x"4E", x"4E", x"4E", x"4D", x"92", x"DB", x"DB", x"DB", x"92", x"6D", x"92", x"92", x"92", x"6D", x"B6", x"DB", x"DB", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"68", x"8C", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"8C", x"88", x"B6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"2E", x"4E", x"92", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"68", x"B6", x"DB", x"B6", x"92", x"92", x"24", x"00", x"24", x"24", x"00", x"00", x"24", x"29", x"92", x"B7", x"6E", x"6E", x"6D", x"6E", x"B6", x"B6", x"DB", x"8D", x"91", x"DB", x"8C", x"68", x"68", x"B2", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"B6", x"88", x"68", x"48", x"6D", x"91", x"B6", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"92", x"DB", x"DB", x"DB", x"B6", x"92", x"92", x"DB", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"91", x"8D", x"B1", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"B1", x"91", x"D6", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"2E", x"4E", x"92", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"88", x"B6", x"DB", x"B6", x"92", x"92", x"6E", x"25", x"29", x"29", x"25", x"25", x"29", x"49", x"92", x"DB", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"DB", x"B6", x"B6", x"DB", x"8C", x"88", x"68", x"B6", x"DA", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"B6", x"DB", x"DB", x"B6", x"92", x"92", x"92", x"92", x"92", x"6D", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"2E", x"4E", x"92", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"68", x"88", x"88", x"8C", x"B6", x"DB", x"B6", x"91", x"6D", x"69", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"92", x"B6", x"6D", x"6D", x"92", x"B6", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"8C", x"68", x"68", x"91", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B6", x"B1", x"88", x"68", x"68", x"6D", x"91", x"B6", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"49", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"96", x"DB", x"DB", x"B6", x"92", x"92", x"B6", x"DB", x"B6", x"B6", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"2E", x"4E", x"96", x"88", x"88", x"88", x"88", x"88", x"68", x"44", x"44", x"44", x"44", x"44", x"68", x"88", x"8D", x"B6", x"DB", x"B6", x"92", x"6D", x"44", x"44", x"44", x"44", x"44", x"44", x"48", x"92", x"B6", x"49", x"6E", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"BB", x"DB", x"8C", x"88", x"68", x"68", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"B7", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"29", x"29", x"29", x"2E", x"4E", x"4E", x"6E", x"92", x"B6", x"DB", x"B6", x"92", x"92", x"6D", x"92", x"92", x"92", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"25", x"2E", x"4F", x"4F", x"4F", x"2E", x"2E", x"2E", x"4E", x"72", x"8D", x"8C", x"88", x"88", x"88", x"88", x"68", x"68", x"44", x"44", x"44", x"44", x"44", x"44", x"68", x"B2", x"D6", x"D6", x"B6", x"92", x"91", x"91", x"91", x"91", x"91", x"91", x"B6", x"B6", x"6D", x"69", x"6D", x"8D", x"92", x"B2", x"B6", x"B6", x"D6", x"B6", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"68", x"68", x"6D", x"8D", x"B6", x"48", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"92", x"B6", x"DB", x"B6", x"B6", x"92", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"49", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"29", x"2A", x"2E", x"4F", x"4F", x"2F", x"2E", x"4E", x"4E", x"2E", x"4E", x"6E", x"6D", x"8C", x"8D", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8C", x"8D", x"91", x"8D", x"8D", x"91", x"91", x"91", x"91", x"91", x"91", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"91", x"91", x"B1", x"B1", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8C", x"68", x"6D", x"92", x"92", x"48", x"68", x"B6", x"B6", x"49", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"4E", x"4E", x"4E", x"72", x"B6", x"DB", x"DB", x"B6", x"92", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"B6", x"6D", x"24", x"00", x"24", x"24", x"24", x"24", x"24", x"49", x"92", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"6D", x"49", x"2A", x"2A", x"2A", x"2A", x"2A", x"2A", x"2A", x"2A", x"2A", x"4A", x"6E", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"B2", x"91", x"6D", x"92", x"91", x"68", x"68", x"68", x"B6", x"DB", x"6D", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"B6", x"DB", x"DB", x"B6", x"92", x"B6", x"92", x"92", x"92", x"6D", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"24", x"49", x"6D", x"6D", x"6D", x"49", x"49", x"6D", x"6D", x"92", x"6D", x"92", x"92", x"92", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"6D", x"6D", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"91", x"92", x"91", x"8D", x"6D", x"8D", x"6D", x"91", x"6D", x"6D", x"68", x"68", x"68", x"68", x"68", x"88", x"B2", x"92", x"49", x"68", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"25", x"29", x"29", x"4E", x"4E", x"4E", x"72", x"96", x"DB", x"DB", x"B6", x"92", x"92", x"B6", x"DB", x"B6", x"B6", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"6D", x"6D", x"92", x"92", x"B6", x"92", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"B2", x"B6", x"B6", x"D6", x"B6", x"D6", x"92", x"49", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"B6", x"8D", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"8C", x"8D", x"92", x"6D", x"68", x"68", x"64", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"29", x"29", x"29", x"2E", x"4E", x"4E", x"6E", x"92", x"B6", x"DB", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"92", x"B6", x"92", x"92", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"B6", x"92", x"92", x"92", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"92", x"B6", x"92", x"B6", x"B6", x"B6", x"B6", x"92", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"8D", x"91", x"B1", x"B1", x"B1", x"B1", x"B1", x"91", x"8D", x"92", x"B6", x"DB", x"DB", x"DB", x"DB", x"B6", x"B1", x"B1", x"91", x"91", x"91", x"91", x"91", x"91", x"8D", x"8D", x"8D", x"B1", x"B2", x"92", x"6D", x"48", x"68", x"68", x"6C", x"48", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"29", x"25", x"29", x"2E", x"2E", x"4E", x"4E", x"92", x"B6", x"DB", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"B6", x"92", x"92", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"92", x"92", x"B6", x"92", x"92", x"B6", x"92", x"B6", x"B6", x"92", x"B6", x"B6", x"B6", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"8D", x"68", x"6C", x"68", x"6C", x"68", x"68", x"68", x"68", x"6C", x"6D", x"6D", x"48", x"24"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"24", x"24", x"24", x"24", x"49", x"49", x"25", x"25", x"25", x"29", x"29", x"49", x"4D", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"8D", x"49", x"48", x"48", x"48", x"48", x"49", x"48", x"49", x"48", x"69", x"48", x"69", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"91", x"8D", x"68", x"48", x"FF", x"48", x"44"),
(x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"48", x"48", x"48", x"48", x"48", x"48", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6C", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6C", x"44", x"92", x"48", x"44", x"00", x"00")
);

-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (
("000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;
  end process;
end behav;		

--generated with PNGtoVHDL tool by Ben Wellingstein
